../riscv.ckt