NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.00025 ;

DIVIDERCHAR "/" ;



LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 0.036 ;
  WIDTH 0.018 ;
  AREA 0.00067 ;
  SPACING 0.018 ;
  SPACING 0.018 RANGE 0.018 1.00 ;
  SPACING 0.105 RANGE 1.00 2.50 ;
  SPACING 0.185 RANGE 2.50 25000 ;
END M1

LAYER V1
  TYPE CUT ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.036 0.036 ;
  WIDTH 0.018 ;
  AREA 0.00067 ;
  MINSIZE 0.037 0.018 ; 
  SPACING 0.018 ;
  SPACING 0.018 RANGE 0.018 1.00 ;
  SPACING 0.105 RANGE 1.00 2.50 ;
  SPACING 0.185 RANGE 2.50 25000 ;
END M2

LAYER V2
  TYPE CUT ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.054 0.036 ;
  WIDTH 0.018 ;
  AREA 0.00067 ;
  SPACING 0.036 ;
  SPACING 0.036 RANGE 0.036 1.00 ;
  SPACING 0.105 RANGE 1.00 2.50 ;
  SPACING 0.185 RANGE 2.50 25000 ;
END M3

LAYER V3
  TYPE CUT ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.048 0.048 ;
  WIDTH 0.024 ;
  AREA 0.002 ;
  SPACING 0.024 ;
  SPACING 0.024 RANGE 0.024 1.00 ;
  SPACING 0.05 RANGE 1.00 2.50 ;
  SPACING 0.105 RANGE 2.50 6.25 ;
  SPACING 0.185 RANGE 6.25 25000 ;
END M4

LAYER V4
  TYPE CUT ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.048 0.048 ;
  WIDTH 0.024 ;
  AREA 0.002 ;
  SPACING 0.024 ;
  SPACING 0.024 RANGE 0.024 1.00 ;
  SPACING 0.05 RANGE 1.00 2.50 ;
  SPACING 0.105 RANGE 2.50 6.25 ;
  SPACING 0.185 RANGE 6.25 25000 ;
END M5

LAYER V5
  TYPE CUT ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 0.064 ;
  WIDTH 0.032 ;
  AREA 0.0021875 ;
  SPACING 0.032 ;
  SPACING 0.032 RANGE 0.032 1.00 ;
  SPACING 0.05 RANGE 1.00 2.00 ;
  SPACING 0.105 RANGE 2.00 6.25 ;
  SPACING 0.185 RANGE 6.25 25000 ;
  END M6


LAYER V6
  TYPE CUT ;
END V6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 0.064 ;
  WIDTH 0.032 ;
  AREA 0.0021875 ;
  SPACING 0.032 ;
  SPACING 0.032 RANGE 0.032 1.00 ;
  SPACING 0.05 RANGE 1.00 2.00 ;
  SPACING 0.105 RANGE 2.00 6.25 ;
  SPACING 0.185 RANGE 6.25 25000 ;
  END M7

LAYER V7
  TYPE CUT ;
END V7

LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 0.08 ;
  WIDTH 0.04 ;
  AREA 0.0025 ;  
  SPACING 0.04 ;
  SPACING 0.04 RANGE 0.04 1.00 ;
  SPACING 0.0625 RANGE 1.00 2.00 ;
  SPACING 0.125 RANGE 2.00 6.25 ;
  SPACING 0.2 RANGE 6.25 25000 ;
  END M8

LAYER V8
  TYPE CUT ;
END V8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 0.08 ;
  WIDTH 0.04 ;
  AREA 0.0025 ;  
  SPACING 0.04 ;
  SPACING 0.04 RANGE 0.04 1.00 ;
  SPACING 0.0625 RANGE 1.00 2.00 ;
  SPACING 0.125 RANGE 2.00 6.25 ;
  SPACING 0.2 RANGE 6.25 25000 ;
  END M9

LAYER V9
  TYPE CUT ;
END V9


LAYER Pad
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 0.08 ;
  WIDTH 0.04 ;
  SPACING 0.04 ;
END Pad



LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

SPACING
  SAMENET M1  M1    0.025 STACK ;
  SAMENET M2  M2    0.04 STACK ;
  SAMENET M3  M3    0.04 STACK ;
  SAMENET M4  M4    0.0625 STACK ;
  SAMENET M5  M5    0.0625 STACK ;
  SAMENET M6  M6    0.1 STACK ;
  SAMENET M7  M7    0.1 STACK ;
  SAMENET M8  M8    0.125 STACK ;
  SAMENET M9  M9    0.125 STACK ;
  SAMENET V1  V1    0.018 ;
  SAMENET V2  V2    0.018 ;
  SAMENET V3  V3    0.018 ;
  SAMENET V4  V4    0.034 ;
  SAMENET V5  V5    0.034 ;
  SAMENET V6  V6    0.046 ;
  SAMENET V7  V7    0.046 ;
  SAMENET V8  V8    0.057 ;
  SAMENET V9  V9    0.057 ;
  SAMENET V1  V2    0.00 STACK ;
  SAMENET V2  V3    0.00 STACK ;
  SAMENET V3  V4    0.00 STACK ;
  SAMENET V4  V5    0.00 STACK ;
  SAMENET V5  V6    0.00 STACK ;
  SAMENET V6  V7    0.00 STACK ;
  SAMENET V7  V8    0.00 STACK ;
  SAMENET V8  V9    0.00 STACK ;
  SAMENET V1  V3    0.00 STACK ;
  SAMENET V2  V4    0.00 STACK ;
  SAMENET V3  V5    0.00 STACK ;
  SAMENET V4  V6    0.00 STACK ;
  SAMENET V5  V7    0.00 STACK ;
  SAMENET V6  V8    0.00 STACK ;
  SAMENET V7  V9    0.00 STACK ;
  SAMENET V1  V4    0.00 STACK ;
  SAMENET V2  V5    0.00 STACK ;
  SAMENET V3  V6    0.00 STACK ;
  SAMENET V4  V7    0.00 STACK ;
  SAMENET V5  V8    0.00 STACK ;
  SAMENET V6  V9    0.00 STACK ;
  SAMENET V1  V5    0.00 STACK ;
  SAMENET V2  V6    0.00 STACK ;
  SAMENET V3  V7    0.00 STACK ;
  SAMENET V4  V8    0.00 STACK ;
  SAMENET V5  V9    0.00 STACK ;
  SAMENET V1  V6    0.00 STACK ;
  SAMENET V2  V7    0.00 STACK ;
  SAMENET V3  V8    0.00 STACK ;
  SAMENET V4  V9    0.00 STACK ;
  SAMENET V1  V7    0.00 STACK ;
  SAMENET V2  V8    0.00 STACK ;
  SAMENET V3  V9    0.00 STACK ;
  SAMENET V1  V8    0.00 STACK ;
  SAMENET V2  V9    0.00 STACK ;
  SAMENET V1  V8    0.00 STACK ;
END SPACING


VIA via9 DEFAULT
  LAYER M9 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER V9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER Pad  ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
END via9

VIA via8 DEFAULT
  LAYER M8 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER V8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER M9 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
END via8

VIA via7 DEFAULT
  LAYER M7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER V7 ;
    RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
END via7

VIA via6 DEFAULT
  LAYER M6 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER V6 ;
    RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M7 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END via6

VIA via5 DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER V5 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER M6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
END via5

VIA via4 DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER V4 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER M5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
END via4

VIA via3 DEFAULT
  LAYER M4 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER V3 ;
    RECT -0.036 -0.036 0.036 0.036 ;
  LAYER M3 ;
    RECT -0.06 -0.06 0.06 0.06 ;
END via3

VIA via2 DEFAULT
  LAYER M3 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER V2 ;
    RECT -0.009 -0.009 0.009 0.009 ; 
  LAYER M2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
END via2

VIA via1 DEFAULT
  LAYER M1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER V1 ;
    RECT -0.009 -0.009 0.009 0.009 ;  
END via1


VIARULE via1Array GENERATE
  LAYER M1 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.01125 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION HORIZONTAL ;
    OVERHANG 0.01125 ;
    METALOVERHANG 0 ;
  LAYER V1 ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.018 BY 0.018 ;
END via1Array

VIARULE via2Array GENERATE
  LAYER M3 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION HORIZONTAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER V2 ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.018 BY 0.018 ;
END via2Array

VIARULE via3Array GENERATE
  LAYER M3 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER V3 ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.018 BY 0.018 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER M5 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER V4 ;
    RECT -0.012 -0.012 0.012 0.012 ;
    SPACING 0.034 BY 0.034 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER M5 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01125 ;
    METALOVERHANG 0 ;
  LAYER V5 ;
    RECT -0.012 -0.012 0.012 0.012 ;
    SPACING 0.034 BY 0.034 ;
END via5Array

VIARULE via6Array GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER M7 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.01125 ;
    METALOVERHANG 0 ;
  LAYER V6 ;
    RECT -0.0016 -0.0016 0.0016 0.0016 ;
    SPACING 0.046 BY 0.046 ;
END via6Array

VIARULE via7Array GENERATE
  LAYER M7 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER M8 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01125 ;
    METALOVERHANG 0 ;
  LAYER V7 ;
    RECT -0.0016 -0.0016 0.0016 0.0016 ;
    SPACING 0.046 BY 0.046 ;
END via7Array

VIARULE via8Array GENERATE
  LAYER M8 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER M9 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.01125 ;
    METALOVERHANG 0 ;
  LAYER V8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
    SPACING 0.057 BY 0.057 ;
END via8Array

VIARULE via9Array GENERATE
  LAYER M9 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.0075 ;
    METALOVERHANG 0 ;
  LAYER Pad ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01125 ;
    METALOVERHANG 0 ;
  LAYER V9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
    SPACING 0.057 BY 0.057 ;
END via9Array

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION VERTICAL ;
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION VERTICAL ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER M5 ;
    DIRECTION VERTICAL ;
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
END TURNM6

VIARULE TURNM7 GENERATE
  LAYER M7 ;
    DIRECTION VERTICAL ;
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
END TURNM7

VIARULE TURNM8 GENERATE
  LAYER M8 ;
    DIRECTION HORIZONTAL ;
  LAYER M8 ;
    DIRECTION VERTICAL ;
END TURNM8

VIARULE TURNM9 GENERATE
  LAYER M9 ;
    DIRECTION VERTICAL ;
  LAYER M9 ;
    DIRECTION HORIZONTAL ;
END TURNM9

VIARULE TURNPad GENERATE
  LAYER Pad ;
    DIRECTION HORIZONTAL ;
  LAYER Pad ;
    DIRECTION VERTICAL ;
END TURNPad


SITE  coreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.036 BY 0.288 ;
END  coreSite



MACRO AOAI211_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211_1x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.333 0 0.351 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.33 0.27 0.348 0.288 ;
        RECT 0.366 0.27 0.384 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.085 0.171 0.103 ;
        RECT 0.018 0.189 0.117 0.207 ;
        RECT 0.018 0.085 0.036 0.207 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.099 0.037 0.279 0.055 ;
      RECT 0.153 0.233 0.279 0.251 ;
  END
END AOAI211_1x

MACRO AOAI211_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211_2x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.214 0 0.232 0.018 ;
        RECT 0.337 0 0.355 0.018 ;
        RECT 0.577 0 0.595 0.018 ;
        RECT 0.621 0 0.639 0.018 ;
        RECT 0.657 0 0.675 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.054 0.27 0.072 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.5275 0.27 0.5455 0.288 ;
        RECT 0.6175 0.27 0.6355 0.288 ;
        RECT 0.654 0.27 0.672 0.288 ;
        RECT 0.69 0.27 0.708 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.32 0.036 0.441 0.054 ;
        RECT 0.018 0.0795 0.338 0.0975 ;
        RECT 0.32 0.036 0.338 0.0975 ;
        RECT 0.018 0.198 0.279 0.216 ;
        RECT 0.018 0.0795 0.036 0.216 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.369 0.082 0.601 0.1 ;
      RECT 0.5215 0.036 0.558 0.054 ;
      RECT 0.207 0.234 0.549 0.252 ;
      RECT 0.2515 0.036 0.288 0.054 ;
      RECT 0.1435 0.036 0.18 0.054 ;
      RECT 0.045 0.036 0.0815 0.054 ;
    LAYER M2 ;
      RECT 0.047 0.036 0.547 0.054 ;
    LAYER V1 ;
      RECT 0.529 0.036 0.547 0.054 ;
      RECT 0.268 0.036 0.286 0.054 ;
      RECT 0.16 0.036 0.178 0.054 ;
      RECT 0.047 0.036 0.065 0.054 ;
  END
END AOAI211_2x

MACRO AOAI211_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211_3x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.268 0 0.286 0.018 ;
        RECT 0.391 0 0.409 0.018 ;
        RECT 0.729 0 0.747 0.018 ;
        RECT 0.765 0 0.783 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.054 0.27 0.072 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.455 0.27 0.473 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.7255 0.27 0.7435 0.288 ;
        RECT 0.762 0.27 0.78 0.288 ;
        RECT 0.798 0.27 0.816 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.128 0.576 0.158 ;
      LAYER M2 ;
        RECT 0.558 0.125 0.576 0.158 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.046 0.495 0.064 ;
        RECT 0.018 0.1875 0.333 0.2055 ;
        RECT 0.018 0.046 0.036 0.2055 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.526 0.046 0.711 0.064 ;
      RECT 0.261 0.234 0.711 0.252 ;
      RECT 0.423 0.082 0.657 0.1 ;
      RECT 0.099 0.082 0.333 0.1 ;
    LAYER M2 ;
      RECT 0.2775 0.082 0.333 0.1 ;
      RECT 0.315 0.046 0.333 0.1 ;
      RECT 0.315 0.046 0.546 0.064 ;
    LAYER V1 ;
      RECT 0.528 0.046 0.546 0.064 ;
      RECT 0.2775 0.082 0.2955 0.1 ;
  END
END AOAI211_3x

MACRO AOAI211_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211_5x 0 0 ;
  SIZE 1.296 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.296 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.296 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.376 0 0.394 0.018 ;
        RECT 0.607 0 0.625 0.018 ;
        RECT 1.161 0 1.179 0.018 ;
        RECT 1.197 0 1.215 0.018 ;
        RECT 1.273 0 1.291 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.054 0.27 0.072 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.671 0.27 0.689 0.288 ;
        RECT 0.9055 0.27 0.9235 0.288 ;
        RECT 1.1575 0.27 1.1755 0.288 ;
        RECT 1.194 0.27 1.212 0.288 ;
        RECT 1.23 0.27 1.248 0.288 ;
        RECT 1.273 0.27 1.291 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.882 0.128 0.9 0.158 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.046 0.819 0.064 ;
        RECT 0.018 0.1875 0.549 0.2055 ;
        RECT 0.018 0.046 0.036 0.2055 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.85 0.046 1.143 0.064 ;
      RECT 0.369 0.234 1.143 0.252 ;
      RECT 0.639 0.082 1.089 0.1 ;
      RECT 0.099 0.082 0.549 0.1 ;
    LAYER M2 ;
      RECT 0.4935 0.082 0.549 0.1 ;
      RECT 0.531 0.046 0.549 0.1 ;
      RECT 0.531 0.046 0.87 0.064 ;
    LAYER V1 ;
      RECT 0.852 0.046 0.87 0.064 ;
      RECT 0.4935 0.082 0.5115 0.1 ;
  END
END AOAI211_5x

MACRO AOAI211_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211_7x 0 0 ;
  SIZE 1.728 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.728 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.728 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.484 0 0.502 0.018 ;
        RECT 0.793 0 0.811 0.018 ;
        RECT 1.593 0 1.611 0.018 ;
        RECT 1.629 0 1.647 0.018 ;
        RECT 1.705 0 1.723 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.054 0.27 0.072 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.527 0.27 0.545 0.288 ;
        RECT 0.887 0.27 0.905 0.288 ;
        RECT 1.2295 0.27 1.2475 0.288 ;
        RECT 1.5895 0.27 1.6075 0.288 ;
        RECT 1.626 0.27 1.644 0.288 ;
        RECT 1.662 0.27 1.68 0.288 ;
        RECT 1.705 0.27 1.723 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.128 1.224 0.158 ;
      LAYER M2 ;
        RECT 1.206 0.125 1.224 0.158 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.046 1.143 0.064 ;
        RECT 0.018 0.1875 0.765 0.2055 ;
        RECT 0.018 0.046 0.036 0.2055 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 1.174 0.046 1.575 0.064 ;
      RECT 0.477 0.234 1.575 0.252 ;
      RECT 0.855 0.082 1.521 0.1 ;
      RECT 0.099 0.082 0.765 0.1 ;
    LAYER M2 ;
      RECT 0.7095 0.082 0.765 0.1 ;
      RECT 0.747 0.046 0.765 0.1 ;
      RECT 0.747 0.046 1.194 0.064 ;
    LAYER V1 ;
      RECT 1.176 0.046 1.194 0.064 ;
      RECT 0.7095 0.082 0.7275 0.1 ;
  END
END AOAI211_7x

MACRO AOI21_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_1x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.351 0 0.369 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.3475 0.27 0.3655 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.229 0.252 0.247 ;
        RECT 0.234 0.041 0.252 0.247 ;
        RECT 0.045 0.041 0.252 0.059 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.171 0.247 ;
  END
END AOI21_1x

MACRO AOI21_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_2x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.177 0 0.195 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.567 0 0.585 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.5635 0.27 0.5815 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.1835 0.522 0.2015 ;
        RECT 0.504 0.085 0.522 0.2015 ;
        RECT 0.099 0.085 0.522 0.103 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.099 0.229 0.495 0.247 ;
      RECT 0.045 0.041 0.279 0.059 ;
  END
END AOI21_2x

MACRO AOI21_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_3x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.231 0 0.249 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.675 0 0.693 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.6715 0.27 0.6895 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.1835 0.576 0.2015 ;
        RECT 0.558 0.085 0.576 0.2015 ;
        RECT 0.045 0.085 0.576 0.103 ;
      LAYER M2 ;
        RECT 0.558 0.125 0.576 0.158 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.495 0.247 ;
      RECT 0.099 0.041 0.333 0.059 ;
  END
END AOI21_3x

MACRO AOI21_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_5x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.339 0 0.357 0.018 ;
        RECT 0.619 0 0.637 0.018 ;
        RECT 0.999 0 1.017 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.617 0.27 0.635 0.288 ;
        RECT 0.9955 0.27 1.0135 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.639 0.1835 0.9 0.2015 ;
        RECT 0.882 0.085 0.9 0.2015 ;
        RECT 0.045 0.085 0.9 0.103 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.819 0.247 ;
      RECT 0.099 0.041 0.549 0.059 ;
  END
END AOI21_5x

MACRO AOI21_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_7x 0 0 ;
  SIZE 1.404 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.404 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.404 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.447 0 0.465 0.018 ;
        RECT 0.835 0 0.853 0.018 ;
        RECT 1.323 0 1.341 0.018 ;
        RECT 1.381 0 1.399 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.404 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.404 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.833 0.27 0.851 0.288 ;
        RECT 1.3195 0.27 1.3375 0.288 ;
        RECT 1.381 0.27 1.399 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.1835 1.224 0.2015 ;
        RECT 1.206 0.085 1.224 0.2015 ;
        RECT 0.045 0.085 1.224 0.103 ;
      LAYER M2 ;
        RECT 1.206 0.125 1.224 0.158 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 1.143 0.247 ;
      RECT 0.099 0.041 0.765 0.059 ;
  END
END AOI21_7x

MACRO AOI22_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_1x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.348 0 0.366 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.3415 0.27 0.3595 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.189 0.306 0.207 ;
        RECT 0.288 0.041 0.306 0.207 ;
        RECT 0.045 0.041 0.306 0.059 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.233 0.279 0.251 ;
  END
END AOI22_1x

MACRO AOI22_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_2x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.256 0 0.274 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.531 0 0.549 0.018 ;
        RECT 0.621 0 0.639 0.018 ;
        RECT 0.672 0 0.69 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.5275 0.27 0.5455 0.288 ;
        RECT 0.6175 0.27 0.6355 0.288 ;
        RECT 0.6655 0.27 0.6835 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.369 0.189 0.63 0.207 ;
        RECT 0.612 0.085 0.63 0.207 ;
        RECT 0.099 0.085 0.63 0.103 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.369 0.049 0.603 0.067 ;
      RECT 0.099 0.233 0.549 0.251 ;
      RECT 0.045 0.049 0.279 0.067 ;
  END
END AOI22_2x

MACRO AOI22_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_3x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.729 0 0.747 0.018 ;
        RECT 0.78 0 0.798 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.7255 0.27 0.7435 0.288 ;
        RECT 0.7735 0.27 0.7915 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.128 0.576 0.158 ;
      LAYER M2 ;
        RECT 0.558 0.125 0.576 0.158 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.189 0.738 0.207 ;
        RECT 0.72 0.085 0.738 0.207 ;
        RECT 0.045 0.085 0.738 0.103 ;
      LAYER M2 ;
        RECT 0.72 0.125 0.738 0.158 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.233 0.711 0.251 ;
      RECT 0.423 0.049 0.657 0.067 ;
      RECT 0.099 0.049 0.333 0.067 ;
  END
END AOI22_3x

MACRO AOI22_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_5x 0 0 ;
  SIZE 1.296 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.296 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.296 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.619 0 0.637 0.018 ;
        RECT 0.909 0 0.927 0.018 ;
        RECT 1.161 0 1.179 0.018 ;
        RECT 1.212 0 1.23 0.018 ;
        RECT 1.273 0 1.291 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.617 0.27 0.635 0.288 ;
        RECT 0.9055 0.27 0.9235 0.288 ;
        RECT 1.1575 0.27 1.1755 0.288 ;
        RECT 1.2055 0.27 1.2235 0.288 ;
        RECT 1.273 0.27 1.291 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.882 0.128 0.9 0.158 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.639 0.189 1.17 0.207 ;
        RECT 1.152 0.085 1.17 0.207 ;
        RECT 0.045 0.085 1.17 0.103 ;
      LAYER M2 ;
        RECT 1.152 0.125 1.17 0.158 ;
      LAYER M3 ;
        RECT 1.152 0.126 1.17 0.158 ;
      LAYER V1 ;
        RECT 1.152 0.13 1.17 0.148 ;
      LAYER V2 ;
        RECT 1.152 0.135 1.17 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.233 1.143 0.251 ;
      RECT 0.639 0.049 1.089 0.067 ;
      RECT 0.099 0.049 0.549 0.067 ;
  END
END AOI22_5x

MACRO AOI22_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_7x 0 0 ;
  SIZE 1.728 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.728 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.728 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.835 0 0.853 0.018 ;
        RECT 1.233 0 1.251 0.018 ;
        RECT 1.593 0 1.611 0.018 ;
        RECT 1.644 0 1.662 0.018 ;
        RECT 1.705 0 1.723 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.833 0.27 0.851 0.288 ;
        RECT 1.2295 0.27 1.2475 0.288 ;
        RECT 1.5895 0.27 1.6075 0.288 ;
        RECT 1.6375 0.27 1.6555 0.288 ;
        RECT 1.705 0.27 1.723 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.128 1.224 0.158 ;
      LAYER M2 ;
        RECT 1.206 0.125 1.224 0.158 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.189 1.602 0.207 ;
        RECT 1.584 0.085 1.602 0.207 ;
        RECT 0.045 0.085 1.602 0.103 ;
      LAYER M2 ;
        RECT 1.584 0.125 1.602 0.158 ;
      LAYER M3 ;
        RECT 1.584 0.126 1.602 0.158 ;
      LAYER V1 ;
        RECT 1.584 0.13 1.602 0.148 ;
      LAYER V2 ;
        RECT 1.584 0.135 1.602 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.233 1.575 0.251 ;
      RECT 0.855 0.049 1.521 0.067 ;
      RECT 0.099 0.049 0.765 0.067 ;
  END
END AOI22_7x

MACRO BUFF_12x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_12x 0 0 ;
  SIZE 1.512 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.512 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.512 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.3655 0 0.3835 0.018 ;
        RECT 0.4735 0 0.4915 0.018 ;
        RECT 0.5815 0 0.5995 0.018 ;
        RECT 0.709 0 0.727 0.018 ;
        RECT 0.799 0 0.817 0.018 ;
        RECT 0.907 0 0.925 0.018 ;
        RECT 1.015 0 1.033 0.018 ;
        RECT 1.123 0 1.141 0.018 ;
        RECT 1.231 0 1.249 0.018 ;
        RECT 1.339 0 1.357 0.018 ;
        RECT 1.375 0 1.393 0.018 ;
        RECT 1.4125 0 1.4305 0.018 ;
        RECT 1.449 0 1.467 0.018 ;
        RECT 1.489 0 1.507 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.512 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.512 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.707 0.27 0.725 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.229 0.27 1.247 0.288 ;
        RECT 1.337 0.27 1.355 0.288 ;
        RECT 1.373 0.27 1.391 0.288 ;
        RECT 1.409 0.27 1.427 0.288 ;
        RECT 1.4455 0.27 1.4635 0.288 ;
        RECT 1.489 0.27 1.507 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.747 0.229 1.386 0.247 ;
        RECT 1.368 0.041 1.386 0.247 ;
        RECT 0.747 0.041 1.386 0.059 ;
      LAYER M2 ;
        RECT 1.368 0.125 1.386 0.158 ;
      LAYER M3 ;
        RECT 1.368 0.126 1.386 0.158 ;
      LAYER V1 ;
        RECT 1.368 0.13 1.386 0.148 ;
      LAYER V2 ;
        RECT 1.368 0.135 1.386 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.657 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.72 0.085 0.738 0.153 ;
      RECT 0.018 0.085 0.738 0.103 ;
  END
END BUFF_12x

MACRO BUFF_16x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_16x 0 0 ;
  SIZE 1.944 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.944 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.944 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.3655 0 0.3835 0.018 ;
        RECT 0.4735 0 0.4915 0.018 ;
        RECT 0.5815 0 0.5995 0.018 ;
        RECT 0.6895 0 0.7075 0.018 ;
        RECT 0.7975 0 0.8155 0.018 ;
        RECT 0.925 0 0.943 0.018 ;
        RECT 1.015 0 1.033 0.018 ;
        RECT 1.123 0 1.141 0.018 ;
        RECT 1.231 0 1.249 0.018 ;
        RECT 1.339 0 1.357 0.018 ;
        RECT 1.447 0 1.465 0.018 ;
        RECT 1.555 0 1.573 0.018 ;
        RECT 1.663 0 1.681 0.018 ;
        RECT 1.771 0 1.789 0.018 ;
        RECT 1.807 0 1.825 0.018 ;
        RECT 1.8445 0 1.8625 0.018 ;
        RECT 1.881 0 1.899 0.018 ;
        RECT 1.921 0 1.939 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.944 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.944 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.923 0.27 0.941 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.229 0.27 1.247 0.288 ;
        RECT 1.337 0.27 1.355 0.288 ;
        RECT 1.445 0.27 1.463 0.288 ;
        RECT 1.553 0.27 1.571 0.288 ;
        RECT 1.661 0.27 1.679 0.288 ;
        RECT 1.769 0.27 1.787 0.288 ;
        RECT 1.805 0.27 1.823 0.288 ;
        RECT 1.841 0.27 1.859 0.288 ;
        RECT 1.8775 0.27 1.8955 0.288 ;
        RECT 1.921 0.27 1.939 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.963 0.229 1.818 0.247 ;
        RECT 1.8 0.041 1.818 0.247 ;
        RECT 0.963 0.041 1.818 0.059 ;
      LAYER M2 ;
        RECT 1.8 0.125 1.818 0.158 ;
      LAYER M3 ;
        RECT 1.8 0.126 1.818 0.158 ;
      LAYER V1 ;
        RECT 1.8 0.13 1.818 0.148 ;
      LAYER V2 ;
        RECT 1.8 0.135 1.818 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.873 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.936 0.085 0.954 0.153 ;
      RECT 0.018 0.085 0.954 0.103 ;
  END
END BUFF_16x

MACRO BUFF_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_1x 0 0 ;
  SIZE 0.324 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.324 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.324 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.301 0 0.319 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.301 0.27 0.319 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.153 0.229 0.198 0.247 ;
        RECT 0.18 0.041 0.198 0.247 ;
        RECT 0.153 0.041 0.198 0.059 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.063 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.126 0.085 0.144 0.153 ;
      RECT 0.018 0.085 0.144 0.103 ;
  END
END BUFF_1x

MACRO BUFF_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_2x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.169 0 0.187 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.295 0 0.313 0.018 ;
        RECT 0.3325 0 0.3505 0.018 ;
        RECT 0.369 0 0.387 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.293 0.27 0.311 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.3655 0.27 0.3835 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.229 0.306 0.247 ;
        RECT 0.288 0.041 0.306 0.247 ;
        RECT 0.207 0.041 0.306 0.059 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.117 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.18 0.085 0.198 0.153 ;
      RECT 0.018 0.085 0.198 0.103 ;
  END
END BUFF_2x

MACRO BUFF_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_3x 0 0 ;
  SIZE 0.54 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.54 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.54 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0955 0 0.1135 0.018 ;
        RECT 0.223 0 0.241 0.018 ;
        RECT 0.313 0 0.331 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.4405 0 0.4585 0.018 ;
        RECT 0.477 0 0.495 0.018 ;
        RECT 0.517 0 0.535 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.4735 0.27 0.4915 0.288 ;
        RECT 0.517 0.27 0.535 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.229 0.414 0.247 ;
        RECT 0.396 0.041 0.414 0.247 ;
        RECT 0.261 0.041 0.414 0.059 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.171 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.234 0.085 0.252 0.153 ;
      RECT 0.018 0.085 0.252 0.103 ;
  END
END BUFF_3x

MACRO BUFF_4x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_4x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.277 0 0.295 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.511 0 0.529 0.018 ;
        RECT 0.5485 0 0.5665 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.275 0.27 0.293 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.509 0.27 0.527 0.288 ;
        RECT 0.545 0.27 0.563 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.315 0.229 0.522 0.247 ;
        RECT 0.504 0.041 0.522 0.247 ;
        RECT 0.315 0.041 0.522 0.059 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.225 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.288 0.085 0.306 0.153 ;
      RECT 0.018 0.085 0.306 0.103 ;
  END
END BUFF_4x

MACRO BUFF_6x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_6x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.385 0 0.403 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.691 0 0.709 0.018 ;
        RECT 0.727 0 0.745 0.018 ;
        RECT 0.7645 0 0.7825 0.018 ;
        RECT 0.801 0 0.819 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.383 0.27 0.401 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.725 0.27 0.743 0.288 ;
        RECT 0.761 0.27 0.779 0.288 ;
        RECT 0.7975 0.27 0.8155 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.229 0.738 0.247 ;
        RECT 0.72 0.041 0.738 0.247 ;
        RECT 0.423 0.041 0.738 0.059 ;
      LAYER M2 ;
        RECT 0.72 0.125 0.738 0.158 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.333 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.396 0.085 0.414 0.153 ;
      RECT 0.018 0.085 0.414 0.103 ;
  END
END BUFF_6x

MACRO BUFF_8x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFF_8x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.3655 0 0.3835 0.018 ;
        RECT 0.493 0 0.511 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.691 0 0.709 0.018 ;
        RECT 0.799 0 0.817 0.018 ;
        RECT 0.907 0 0.925 0.018 ;
        RECT 0.943 0 0.961 0.018 ;
        RECT 0.9805 0 0.9985 0.018 ;
        RECT 1.017 0 1.035 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.491 0.27 0.509 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 0.941 0.27 0.959 0.288 ;
        RECT 0.977 0.27 0.995 0.288 ;
        RECT 1.0135 0.27 1.0315 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.531 0.229 0.954 0.247 ;
        RECT 0.936 0.041 0.954 0.247 ;
        RECT 0.531 0.041 0.954 0.059 ;
      LAYER M2 ;
        RECT 0.936 0.125 0.954 0.158 ;
      LAYER M3 ;
        RECT 0.936 0.126 0.954 0.158 ;
      LAYER V1 ;
        RECT 0.936 0.13 0.954 0.148 ;
      LAYER V2 ;
        RECT 0.936 0.135 0.954 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.441 0.247 ;
      RECT 0.018 0.085 0.036 0.247 ;
      RECT 0.504 0.085 0.522 0.153 ;
      RECT 0.018 0.085 0.522 0.103 ;
  END
END BUFF_8x

MACRO DFF_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF_1x 0 0 ;
  SIZE 1.836 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.836 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.836 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.301 0 0.319 0.018 ;
        RECT 0.3575 0 0.3755 0.018 ;
        RECT 0.3935 0 0.4115 0.018 ;
        RECT 0.4295 0 0.4475 0.018 ;
        RECT 0.4655 0 0.4835 0.018 ;
        RECT 0.5015 0 0.5195 0.018 ;
        RECT 0.5375 0 0.5555 0.018 ;
        RECT 0.5735 0 0.5915 0.018 ;
        RECT 0.61 0 0.628 0.018 ;
        RECT 0.6535 0 0.6715 0.018 ;
        RECT 0.7085 0 0.7265 0.018 ;
        RECT 0.7445 0 0.7625 0.018 ;
        RECT 0.7805 0 0.7985 0.018 ;
        RECT 0.8165 0 0.8345 0.018 ;
        RECT 0.8525 0 0.8705 0.018 ;
        RECT 0.8885 0 0.9065 0.018 ;
        RECT 0.9245 0 0.9425 0.018 ;
        RECT 0.961 0 0.979 0.018 ;
        RECT 1.0045 0 1.0225 0.018 ;
        RECT 1.0635 0 1.0815 0.018 ;
        RECT 1.0995 0 1.1175 0.018 ;
        RECT 1.1355 0 1.1535 0.018 ;
        RECT 1.1715 0 1.1895 0.018 ;
        RECT 1.2075 0 1.2255 0.018 ;
        RECT 1.2435 0 1.2615 0.018 ;
        RECT 1.2795 0 1.2975 0.018 ;
        RECT 1.316 0 1.334 0.018 ;
        RECT 1.3595 0 1.3775 0.018 ;
        RECT 1.409 0 1.427 0.018 ;
        RECT 1.445 0 1.463 0.018 ;
        RECT 1.481 0 1.499 0.018 ;
        RECT 1.517 0 1.535 0.018 ;
        RECT 1.553 0 1.571 0.018 ;
        RECT 1.589 0 1.607 0.018 ;
        RECT 1.625 0 1.643 0.018 ;
        RECT 1.6615 0 1.6795 0.018 ;
        RECT 1.705 0 1.723 0.018 ;
        RECT 1.7595 0 1.7775 0.018 ;
        RECT 1.813 0 1.831 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.836 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.836 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.301 0.27 0.319 0.288 ;
        RECT 0.3575 0.27 0.3755 0.288 ;
        RECT 0.3935 0.27 0.4115 0.288 ;
        RECT 0.4295 0.27 0.4475 0.288 ;
        RECT 0.4655 0.27 0.4835 0.288 ;
        RECT 0.5015 0.27 0.5195 0.288 ;
        RECT 0.5375 0.27 0.5555 0.288 ;
        RECT 0.5735 0.27 0.5915 0.288 ;
        RECT 0.61 0.27 0.628 0.288 ;
        RECT 0.6535 0.27 0.6715 0.288 ;
        RECT 0.7085 0.27 0.7265 0.288 ;
        RECT 0.7445 0.27 0.7625 0.288 ;
        RECT 0.7805 0.27 0.7985 0.288 ;
        RECT 0.8165 0.27 0.8345 0.288 ;
        RECT 0.8525 0.27 0.8705 0.288 ;
        RECT 0.8885 0.27 0.9065 0.288 ;
        RECT 0.9245 0.27 0.9425 0.288 ;
        RECT 0.961 0.27 0.979 0.288 ;
        RECT 1.0045 0.27 1.0225 0.288 ;
        RECT 1.0635 0.27 1.0815 0.288 ;
        RECT 1.0995 0.27 1.1175 0.288 ;
        RECT 1.1355 0.27 1.1535 0.288 ;
        RECT 1.1715 0.27 1.1895 0.288 ;
        RECT 1.2075 0.27 1.2255 0.288 ;
        RECT 1.2435 0.27 1.2615 0.288 ;
        RECT 1.2795 0.27 1.2975 0.288 ;
        RECT 1.316 0.27 1.334 0.288 ;
        RECT 1.3595 0.27 1.3775 0.288 ;
        RECT 1.409 0.27 1.427 0.288 ;
        RECT 1.445 0.27 1.463 0.288 ;
        RECT 1.481 0.27 1.499 0.288 ;
        RECT 1.517 0.27 1.535 0.288 ;
        RECT 1.553 0.27 1.571 0.288 ;
        RECT 1.589 0.27 1.607 0.288 ;
        RECT 1.625 0.27 1.643 0.288 ;
        RECT 1.6615 0.27 1.6795 0.288 ;
        RECT 1.705 0.27 1.723 0.288 ;
        RECT 1.7595 0.27 1.7775 0.288 ;
        RECT 1.813 0.27 1.831 0.288 ;
    END
  END VDD!
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.665 0.228 1.71 0.246 ;
        RECT 1.692 0.039 1.71 0.246 ;
        RECT 1.665 0.039 1.71 0.057 ;
      LAYER M2 ;
        RECT 1.692 0.125 1.71 0.158 ;
      LAYER M3 ;
        RECT 1.692 0.126 1.71 0.158 ;
      LAYER V1 ;
        RECT 1.692 0.13 1.71 0.148 ;
      LAYER V2 ;
        RECT 1.692 0.135 1.71 0.153 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.476 0.123 1.494 0.153 ;
        RECT 0.288 0.128 0.306 0.158 ;
      LAYER M2 ;
        RECT 1.476 0.045 1.494 0.146 ;
        RECT 0.288 0.045 1.494 0.063 ;
        RECT 0.288 0.045 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
        RECT 1.476 0.128 1.494 0.146 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END R
  OBS
    LAYER M1 ;
      RECT 1.503 0.233 1.548 0.251 ;
      RECT 1.53 0.08 1.548 0.251 ;
      RECT 1.368 0.08 1.386 0.153 ;
      RECT 1.368 0.08 1.548 0.098 ;
      RECT 1.26 0.188 1.359 0.206 ;
      RECT 1.26 0.037 1.278 0.206 ;
      RECT 1.179 0.037 1.359 0.055 ;
      RECT 1.098 0.183 1.197 0.201 ;
      RECT 1.098 0.037 1.116 0.201 ;
      RECT 1.017 0.037 1.143 0.055 ;
      RECT 0.963 0.225 1.143 0.243 ;
      RECT 1.044 0.086 1.062 0.243 ;
      RECT 0.963 0.086 1.062 0.104 ;
      RECT 0.831 0.183 1.011 0.201 ;
      RECT 0.99 0.133 1.008 0.201 ;
      RECT 0.639 0.233 0.873 0.251 ;
      RECT 0.774 0.037 0.792 0.251 ;
      RECT 0.693 0.037 0.873 0.055 ;
      RECT 0.585 0.19 0.738 0.208 ;
      RECT 0.72 0.082 0.738 0.208 ;
      RECT 0.639 0.082 0.738 0.1 ;
      RECT 0.423 0.188 0.549 0.206 ;
      RECT 0.45 0.037 0.468 0.206 ;
      RECT 0.423 0.037 0.603 0.055 ;
      RECT 0.342 0.233 0.603 0.251 ;
      RECT 0.342 0.135 0.36 0.251 ;
      RECT 0.153 0.183 0.198 0.201 ;
      RECT 0.18 0.041 0.198 0.201 ;
      RECT 0.369 0.041 0.387 0.102 ;
      RECT 0.153 0.041 0.387 0.059 ;
      RECT 0.234 0.225 0.284 0.243 ;
      RECT 0.234 0.085 0.252 0.243 ;
      RECT 0.234 0.085 0.333 0.103 ;
      RECT 0.018 0.183 0.091 0.201 ;
      RECT 0.018 0.085 0.036 0.201 ;
      RECT 0.126 0.085 0.144 0.153 ;
      RECT 0.018 0.085 0.144 0.103 ;
      RECT 1.638 0.133 1.656 0.163 ;
      RECT 1.422 0.133 1.44 0.163 ;
      RECT 1.314 0.133 1.332 0.163 ;
      RECT 1.179 0.225 1.305 0.243 ;
      RECT 1.152 0.123 1.17 0.153 ;
      RECT 0.936 0.128 0.954 0.156 ;
      RECT 0.882 0.128 0.9 0.156 ;
      RECT 0.666 0.133 0.684 0.163 ;
      RECT 0.612 0.123 0.63 0.153 ;
      RECT 0.558 0.133 0.576 0.163 ;
    LAYER M2 ;
      RECT 1.285 0.225 1.656 0.243 ;
      RECT 1.638 0.14 1.656 0.243 ;
      RECT 1.422 0.14 1.44 0.243 ;
      RECT 0.99 0.183 1.332 0.201 ;
      RECT 1.314 0.14 1.332 0.201 ;
      RECT 1.152 0.082 1.17 0.146 ;
      RECT 0.612 0.082 0.63 0.146 ;
      RECT 0.369 0.082 1.17 0.1 ;
      RECT 0.264 0.225 0.954 0.243 ;
      RECT 0.936 0.136 0.954 0.243 ;
      RECT 0.882 0.136 0.9 0.243 ;
      RECT 0.071 0.183 0.851 0.201 ;
      RECT 0.666 0.14 0.684 0.201 ;
      RECT 0.558 0.14 0.576 0.201 ;
    LAYER V1 ;
      RECT 1.638 0.14 1.656 0.158 ;
      RECT 1.422 0.14 1.44 0.158 ;
      RECT 1.314 0.14 1.332 0.158 ;
      RECT 1.285 0.225 1.303 0.243 ;
      RECT 1.152 0.128 1.17 0.146 ;
      RECT 0.99 0.183 1.008 0.201 ;
      RECT 0.936 0.136 0.954 0.154 ;
      RECT 0.882 0.136 0.9 0.154 ;
      RECT 0.833 0.183 0.851 0.201 ;
      RECT 0.666 0.14 0.684 0.158 ;
      RECT 0.612 0.128 0.63 0.146 ;
      RECT 0.558 0.14 0.576 0.158 ;
      RECT 0.369 0.082 0.387 0.1 ;
      RECT 0.264 0.225 0.282 0.243 ;
      RECT 0.071 0.183 0.089 0.201 ;
  END
END DFF_1x

MACRO FILLER
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER 0 0 ;
  SIZE 0.036 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.036 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.036 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.036 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.036 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
    END
  END VDD!
END FILLER

MACRO INV_12x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_12x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.745 0 0.763 0.018 ;
        RECT 0.781 0 0.799 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.743 0.27 0.761 0.288 ;
        RECT 0.779 0.27 0.797 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.1585 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.2265 0.738 0.2445 ;
        RECT 0.72 0.041 0.738 0.2445 ;
        RECT 0.099 0.041 0.738 0.059 ;
      LAYER M2 ;
        RECT 0.72 0.125 0.738 0.158 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END OUT
END INV_12x

MACRO INV_16x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_16x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.961 0 0.979 0.018 ;
        RECT 0.997 0 1.015 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.959 0.27 0.977 0.288 ;
        RECT 0.995 0.27 1.013 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.1585 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.2265 0.954 0.2445 ;
        RECT 0.936 0.041 0.954 0.2445 ;
        RECT 0.099 0.041 0.954 0.059 ;
      LAYER M2 ;
        RECT 0.936 0.125 0.954 0.158 ;
      LAYER M3 ;
        RECT 0.936 0.126 0.954 0.158 ;
      LAYER V1 ;
        RECT 0.936 0.13 0.954 0.148 ;
      LAYER V2 ;
        RECT 0.936 0.135 0.954 0.153 ;
    END
  END OUT
END INV_16x

MACRO INV_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_1x 0 0 ;
  SIZE 0.324 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.324 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.324 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.241 0 0.259 0.018 ;
        RECT 0.301 0 0.319 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.239 0.27 0.257 0.288 ;
        RECT 0.301 0.27 0.319 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.229 0.144 0.247 ;
        RECT 0.126 0.041 0.144 0.247 ;
        RECT 0.099 0.041 0.144 0.059 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END OUT
END INV_1x

MACRO INV_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_2x 0 0 ;
  SIZE 0.324 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.324 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.324 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.241 0 0.259 0.018 ;
        RECT 0.301 0 0.319 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.239 0.27 0.257 0.288 ;
        RECT 0.301 0.27 0.319 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.2265 0.198 0.2445 ;
        RECT 0.18 0.041 0.198 0.2445 ;
        RECT 0.099 0.041 0.198 0.059 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END OUT
END INV_2x

MACRO INV_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_3x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.349 0 0.367 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.347 0.27 0.365 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.2265 0.252 0.2445 ;
        RECT 0.234 0.041 0.252 0.2445 ;
        RECT 0.099 0.041 0.252 0.059 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END OUT
END INV_3x

MACRO INV_4x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_4x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.313 0 0.331 0.018 ;
        RECT 0.349 0 0.367 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.347 0.27 0.365 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.2265 0.306 0.2445 ;
        RECT 0.288 0.041 0.306 0.2445 ;
        RECT 0.099 0.041 0.306 0.059 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END OUT
END INV_4x

MACRO INV_6x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_6x 0 0 ;
  SIZE 0.54 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.54 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.54 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.421 0 0.439 0.018 ;
        RECT 0.457 0 0.475 0.018 ;
        RECT 0.517 0 0.535 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.455 0.27 0.473 0.288 ;
        RECT 0.517 0.27 0.535 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.2265 0.414 0.2445 ;
        RECT 0.396 0.041 0.414 0.2445 ;
        RECT 0.099 0.041 0.414 0.059 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END OUT
END INV_6x

MACRO INV_8x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_8x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.529 0 0.547 0.018 ;
        RECT 0.565 0 0.583 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.527 0.27 0.545 0.288 ;
        RECT 0.563 0.27 0.581 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.2265 0.522 0.2445 ;
        RECT 0.504 0.041 0.522 0.2445 ;
        RECT 0.099 0.041 0.522 0.059 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END OUT
END INV_8x

MACRO MC_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MC_1x 0 0 ;
  SIZE 0.54 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.54 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.54 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.348 0 0.366 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
        RECT 0.4505 0 0.4685 0.018 ;
        RECT 0.517 0 0.535 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.3415 0.27 0.3595 0.288 ;
        RECT 0.393 0.27 0.411 0.288 ;
        RECT 0.44 0.27 0.458 0.288 ;
        RECT 0.517 0.27 0.535 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.085 0.252 0.153 ;
        RECT 0.126 0.085 0.252 0.103 ;
        RECT 0.126 0.085 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.183 0.306 0.201 ;
        RECT 0.288 0.135 0.306 0.201 ;
        RECT 0.072 0.128 0.09 0.201 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.369 0.225 0.414 0.243 ;
        RECT 0.396 0.041 0.414 0.243 ;
        RECT 0.369 0.041 0.414 0.059 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.342 0.135 0.36 0.165 ;
      RECT 0.207 0.045 0.288 0.063 ;
      RECT 0.207 0.225 0.288 0.243 ;
      RECT 0.045 0.042 0.171 0.06 ;
      RECT 0.045 0.226 0.171 0.244 ;
    LAYER M2 ;
      RECT 0.268 0.225 0.36 0.243 ;
      RECT 0.342 0.045 0.36 0.243 ;
      RECT 0.268 0.045 0.36 0.063 ;
    LAYER V1 ;
      RECT 0.342 0.142 0.36 0.16 ;
      RECT 0.268 0.045 0.286 0.063 ;
      RECT 0.268 0.225 0.286 0.243 ;
  END
END MC_1x

MACRO MC_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MC_2x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.169 0 0.187 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.295 0 0.313 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.621 0 0.639 0.018 ;
        RECT 0.949 0 0.967 0.018 ;
        RECT 0.9905 0 1.0085 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.293 0.27 0.311 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.6175 0.27 0.6355 0.288 ;
        RECT 0.8275 0.27 0.8455 0.288 ;
        RECT 0.933 0.27 0.951 0.288 ;
        RECT 0.98 0.27 0.998 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.123 0.522 0.153 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.082 0.522 0.153 ;
        RECT 0.18 0.082 0.522 0.1 ;
        RECT 0.18 0.082 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
        RECT 0.504 0.128 0.522 0.146 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.135 0.63 0.165 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.183 0.63 0.201 ;
        RECT 0.612 0.135 0.63 0.201 ;
        RECT 0.072 0.125 0.09 0.201 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.612 0.142 0.63 0.16 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.128 0.306 0.158 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.234 0.954 0.252 ;
        RECT 0.936 0.036 0.954 0.252 ;
        RECT 0.855 0.036 0.954 0.054 ;
      LAYER M2 ;
        RECT 0.936 0.125 0.954 0.158 ;
      LAYER M3 ;
        RECT 0.936 0.126 0.954 0.158 ;
      LAYER V1 ;
        RECT 0.936 0.13 0.954 0.148 ;
      LAYER V2 ;
        RECT 0.936 0.135 0.954 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.315 0.19 0.846 0.208 ;
      RECT 0.828 0.08 0.846 0.208 ;
      RECT 0.315 0.08 0.846 0.098 ;
      RECT 0.477 0.044 0.711 0.062 ;
      RECT 0.477 0.226 0.711 0.244 ;
      RECT 0.045 0.044 0.387 0.062 ;
      RECT 0.045 0.226 0.387 0.244 ;
  END
END MC_2x

MACRO MC_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MC_3x 0 0 ;
  SIZE 1.188 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.188 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.188 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.223 0 0.241 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.331 0 0.349 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.693 0 0.711 0.018 ;
        RECT 0.729 0 0.747 0.018 ;
        RECT 0.8815 0 0.8995 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
        RECT 1.0985 0 1.1165 0.018 ;
        RECT 1.165 0 1.183 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.188 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.188 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.6895 0.27 0.7075 0.288 ;
        RECT 0.7255 0.27 0.7435 0.288 ;
        RECT 0.8815 0.27 0.8995 0.288 ;
        RECT 1.041 0.27 1.059 0.288 ;
        RECT 1.088 0.27 1.106 0.288 ;
        RECT 1.165 0.27 1.183 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.123 0.576 0.153 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.558 0.082 0.576 0.153 ;
        RECT 0.234 0.082 0.576 0.1 ;
        RECT 0.234 0.082 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
        RECT 0.558 0.128 0.576 0.146 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.135 0.738 0.165 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.183 0.738 0.201 ;
        RECT 0.72 0.135 0.738 0.201 ;
        RECT 0.072 0.125 0.09 0.201 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.72 0.142 0.738 0.16 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.909 0.226 1.062 0.244 ;
        RECT 1.044 0.039 1.062 0.244 ;
        RECT 0.909 0.039 1.062 0.057 ;
      LAYER M2 ;
        RECT 1.044 0.125 1.062 0.158 ;
      LAYER M3 ;
        RECT 1.044 0.126 1.062 0.158 ;
      LAYER V1 ;
        RECT 1.044 0.13 1.062 0.148 ;
      LAYER V2 ;
        RECT 1.044 0.135 1.062 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.423 0.19 0.9 0.208 ;
      RECT 0.882 0.075 0.9 0.208 ;
      RECT 0.423 0.075 0.9 0.093 ;
      RECT 0.585 0.039 0.819 0.057 ;
      RECT 0.585 0.226 0.819 0.244 ;
      RECT 0.045 0.039 0.495 0.057 ;
      RECT 0.045 0.226 0.495 0.244 ;
  END
END MC_3x

MACRO MC_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MC_5x 0 0 ;
  SIZE 1.836 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.836 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.836 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.331 0 0.349 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.439 0 0.457 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.547 0 0.565 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.619 0 0.637 0.018 ;
        RECT 1.125 0 1.143 0.018 ;
        RECT 1.161 0 1.179 0.018 ;
        RECT 1.4215 0 1.4395 0.018 ;
        RECT 1.705 0 1.723 0.018 ;
        RECT 1.7465 0 1.7645 0.018 ;
        RECT 1.813 0 1.831 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.836 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.836 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.545 0.27 0.563 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.617 0.27 0.635 0.288 ;
        RECT 1.1215 0.27 1.1395 0.288 ;
        RECT 1.1575 0.27 1.1755 0.288 ;
        RECT 1.4215 0.27 1.4395 0.288 ;
        RECT 1.689 0.27 1.707 0.288 ;
        RECT 1.736 0.27 1.754 0.288 ;
        RECT 1.813 0.27 1.831 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.882 0.123 0.9 0.153 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.882 0.082 0.9 0.153 ;
        RECT 0.342 0.082 0.9 0.1 ;
        RECT 0.342 0.082 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
        RECT 0.882 0.128 0.9 0.146 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.135 1.17 0.165 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.183 1.17 0.201 ;
        RECT 1.152 0.135 1.17 0.201 ;
        RECT 0.072 0.125 0.09 0.201 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 1.152 0.142 1.17 0.16 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.449 0.226 1.71 0.244 ;
        RECT 1.692 0.039 1.71 0.244 ;
        RECT 1.449 0.039 1.71 0.057 ;
      LAYER M2 ;
        RECT 1.692 0.125 1.71 0.158 ;
      LAYER M3 ;
        RECT 1.692 0.126 1.71 0.158 ;
      LAYER V1 ;
        RECT 1.692 0.13 1.71 0.148 ;
      LAYER V2 ;
        RECT 1.692 0.135 1.71 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.639 0.19 1.44 0.208 ;
      RECT 1.422 0.075 1.44 0.208 ;
      RECT 0.639 0.075 1.44 0.093 ;
      RECT 0.909 0.039 1.359 0.057 ;
      RECT 0.909 0.226 1.359 0.244 ;
      RECT 0.045 0.039 0.819 0.057 ;
      RECT 0.045 0.226 0.819 0.244 ;
  END
END MC_5x

MACRO MS_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MS_1x 0 0 ;
  SIZE 0.972 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.972 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.972 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.348 0 0.366 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
        RECT 0.4505 0 0.4685 0.018 ;
        RECT 0.61 0 0.628 0.018 ;
        RECT 0.657 0 0.675 0.018 ;
        RECT 0.7275 0 0.7455 0.018 ;
        RECT 0.88 0 0.898 0.018 ;
        RECT 0.949 0 0.967 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.972 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.972 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.3415 0.27 0.3595 0.288 ;
        RECT 0.393 0.27 0.411 0.288 ;
        RECT 0.44 0.27 0.458 0.288 ;
        RECT 0.51 0.27 0.528 0.288 ;
        RECT 0.61 0.27 0.628 0.288 ;
        RECT 0.657 0.27 0.675 0.288 ;
        RECT 0.7275 0.27 0.7455 0.288 ;
        RECT 0.88 0.27 0.898 0.288 ;
        RECT 0.949 0.27 0.967 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.189 0.576 0.207 ;
        RECT 0.558 0.135 0.576 0.207 ;
        RECT 0.342 0.135 0.36 0.207 ;
        RECT 0.234 0.135 0.252 0.165 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.088 0.36 0.155 ;
        RECT 0.234 0.088 0.36 0.106 ;
        RECT 0.126 0.184 0.252 0.202 ;
        RECT 0.234 0.088 0.252 0.202 ;
        RECT 0.126 0.125 0.144 0.202 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
        RECT 0.234 0.137 0.252 0.155 ;
        RECT 0.342 0.137 0.36 0.155 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.135 0.63 0.165 ;
        RECT 0.396 0.13 0.414 0.16 ;
        RECT 0.288 0.135 0.306 0.165 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.225 0.63 0.243 ;
        RECT 0.612 0.137 0.63 0.243 ;
        RECT 0.396 0.137 0.414 0.243 ;
        RECT 0.288 0.137 0.306 0.243 ;
        RECT 0.072 0.125 0.09 0.243 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.288 0.137 0.306 0.155 ;
        RECT 0.396 0.137 0.414 0.155 ;
        RECT 0.612 0.137 0.63 0.155 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.666 0.123 0.684 0.153 ;
        RECT 0.45 0.126 0.468 0.158 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.666 0.052 0.684 0.151 ;
        RECT 0.18 0.052 0.684 0.07 ;
        RECT 0.45 0.052 0.468 0.151 ;
        RECT 0.18 0.052 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
        RECT 0.45 0.133 0.468 0.151 ;
        RECT 0.666 0.133 0.684 0.151 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.747 0.234 0.792 0.252 ;
        RECT 0.774 0.041 0.792 0.252 ;
        RECT 0.747 0.041 0.792 0.059 ;
      LAYER M2 ;
        RECT 0.774 0.125 0.792 0.158 ;
      LAYER M3 ;
        RECT 0.774 0.126 0.792 0.158 ;
      LAYER V1 ;
        RECT 0.774 0.13 0.792 0.148 ;
      LAYER V2 ;
        RECT 0.774 0.135 0.792 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.531 0.2295 0.711 0.2475 ;
      RECT 0.693 0.173 0.711 0.2475 ;
      RECT 0.693 0.173 0.738 0.1915 ;
      RECT 0.72 0.084 0.738 0.1915 ;
      RECT 0.692 0.084 0.738 0.102 ;
      RECT 0.692 0.0385 0.71 0.102 ;
      RECT 0.531 0.0385 0.71 0.0565 ;
      RECT 0.018 0.19 0.225 0.208 ;
      RECT 0.018 0.0815 0.036 0.208 ;
      RECT 0.504 0.0815 0.522 0.153 ;
      RECT 0.018 0.0815 0.522 0.0995 ;
      RECT 0.369 0.0385 0.495 0.0565 ;
      RECT 0.369 0.2295 0.495 0.2475 ;
      RECT 0.045 0.0385 0.171 0.0565 ;
      RECT 0.045 0.2295 0.171 0.2475 ;
  END
END MS_1x

MACRO MS_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MS_2x 0 0 ;
  SIZE 2.052 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 2.052 0.018 ;
      LAYER M2 ;
        RECT 0 0 2.052 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.041 0 0.059 0.018 ;
        RECT 0.167 0 0.185 0.018 ;
        RECT 0.257 0 0.275 0.018 ;
        RECT 0.365 0 0.383 0.018 ;
        RECT 0.491 0 0.5125 0.018 ;
        RECT 0.5815 0 0.603 0.018 ;
        RECT 1.474 0 1.492 0.018 ;
        RECT 1.683 0 1.701 0.018 ;
        RECT 1.96 0 1.978 0.018 ;
        RECT 2.029 0 2.047 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 2.052 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 2.052 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.491 0.27 0.509 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.923 0.27 0.941 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.3395 0.27 1.3575 0.288 ;
        RECT 1.474 0.27 1.492 0.288 ;
        RECT 1.683 0.27 1.701 0.288 ;
        RECT 1.96 0.27 1.978 0.288 ;
        RECT 2.029 0.27 2.047 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.135 1.386 0.163 ;
        RECT 0.828 0.185 1.005 0.203 ;
        RECT 0.828 0.135 0.846 0.203 ;
        RECT 0.504 0.135 0.522 0.165 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.985 0.185 1.386 0.203 ;
        RECT 1.368 0.137 1.386 0.203 ;
        RECT 0.828 0.088 0.846 0.155 ;
        RECT 0.504 0.088 0.846 0.106 ;
        RECT 0.18 0.184 0.522 0.202 ;
        RECT 0.504 0.088 0.522 0.202 ;
        RECT 0.18 0.125 0.198 0.202 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
        RECT 0.504 0.137 0.522 0.155 ;
        RECT 0.828 0.137 0.846 0.155 ;
        RECT 0.985 0.185 1.003 0.203 ;
        RECT 1.368 0.137 1.386 0.155 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.468 0.135 1.499 0.153 ;
        RECT 0.936 0.13 0.954 0.16 ;
        RECT 0.612 0.135 0.63 0.165 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 1.404 0.135 1.494 0.153 ;
        RECT 0.072 0.225 1.422 0.243 ;
        RECT 1.404 0.135 1.422 0.243 ;
        RECT 0.936 0.137 0.954 0.243 ;
        RECT 0.612 0.137 0.63 0.243 ;
        RECT 0.072 0.125 0.09 0.243 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.612 0.137 0.63 0.155 ;
        RECT 0.936 0.137 0.954 0.155 ;
        RECT 1.476 0.135 1.494 0.153 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.1245 1.71 0.153 ;
        RECT 1.044 0.126 1.062 0.158 ;
        RECT 0.288 0.128 0.306 0.158 ;
      LAYER M2 ;
        RECT 1.692 0.045 1.71 0.151 ;
        RECT 0.288 0.045 1.71 0.063 ;
        RECT 1.044 0.045 1.062 0.151 ;
        RECT 0.288 0.045 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
        RECT 1.044 0.133 1.062 0.151 ;
        RECT 1.692 0.133 1.71 0.151 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.827 0.234 1.926 0.252 ;
        RECT 1.908 0.036 1.926 0.252 ;
        RECT 1.827 0.036 1.926 0.054 ;
      LAYER M2 ;
        RECT 1.908 0.125 1.926 0.158 ;
      LAYER M3 ;
        RECT 1.908 0.126 1.926 0.158 ;
      LAYER V1 ;
        RECT 1.908 0.13 1.926 0.148 ;
      LAYER V2 ;
        RECT 1.908 0.135 1.926 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 1.8 0.0815 1.818 0.158 ;
      RECT 1.6135 0.0815 1.818 0.0995 ;
      RECT 1.449 0.091 1.575 0.109 ;
      RECT 1.449 0.045 1.467 0.109 ;
      RECT 1.341 0.045 1.467 0.063 ;
      RECT 0.018 0.19 0.549 0.208 ;
      RECT 0.018 0.0815 0.036 0.208 ;
      RECT 0.018 0.0815 1.1105 0.0995 ;
      RECT 1.503 0.0455 1.737 0.0635 ;
      RECT 1.503 0.1935 1.737 0.2115 ;
      RECT 1.341 0.2295 1.575 0.2475 ;
      RECT 1.179 0.1935 1.472 0.2115 ;
      RECT 1.381 0.0815 1.418 0.0995 ;
      RECT 1.179 0.0815 1.306 0.0995 ;
      RECT 0.801 0.0385 1.251 0.0565 ;
      RECT 0.801 0.2295 1.251 0.2475 ;
      RECT 1.152 0.125 1.17 0.153 ;
      RECT 0.477 0.0405 0.711 0.0585 ;
      RECT 0.477 0.2295 0.711 0.2475 ;
      RECT 0.045 0.0405 0.387 0.0585 ;
      RECT 0.045 0.2295 0.387 0.2475 ;
    LAYER M2 ;
      RECT 1.452 0.1935 1.818 0.2115 ;
      RECT 1.8 0.135 1.818 0.2115 ;
      RECT 1.152 0.0815 1.17 0.151 ;
      RECT 1.0905 0.0815 1.17 0.0995 ;
      RECT 1.286 0.0815 1.6335 0.0995 ;
    LAYER V1 ;
      RECT 1.8 0.135 1.818 0.153 ;
      RECT 1.6155 0.0815 1.6335 0.0995 ;
      RECT 1.452 0.1935 1.47 0.2115 ;
      RECT 1.383 0.0815 1.401 0.0995 ;
      RECT 1.286 0.0815 1.304 0.0995 ;
      RECT 1.152 0.133 1.17 0.151 ;
      RECT 1.0905 0.0815 1.1085 0.0995 ;
  END
END MS_2x

MACRO MS_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MS_3x 0 0 ;
  SIZE 2.376 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 2.376 0.018 ;
      LAYER M2 ;
        RECT 0 0 2.376 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.223 0 0.241 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.888 0 0.906 0.018 ;
        RECT 1.2065 0 1.2245 0.018 ;
        RECT 1.395 0 1.413 0.018 ;
        RECT 1.557 0 1.575 0.018 ;
        RECT 1.69 0 1.708 0.018 ;
        RECT 1.845 0 1.863 0.018 ;
        RECT 2.043 0 2.061 0.018 ;
        RECT 2.284 0 2.302 0.018 ;
        RECT 2.353 0 2.371 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 2.376 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 2.376 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.7435 0.27 0.7615 0.288 ;
        RECT 0.8515 0.27 0.8695 0.288 ;
        RECT 0.9595 0.27 0.9775 0.288 ;
        RECT 1.0675 0.27 1.0855 0.288 ;
        RECT 1.1755 0.27 1.1935 0.288 ;
        RECT 1.2835 0.27 1.3015 0.288 ;
        RECT 1.3375 0.27 1.3555 0.288 ;
        RECT 1.4455 0.27 1.4635 0.288 ;
        RECT 1.5535 0.27 1.5715 0.288 ;
        RECT 1.69 0.27 1.708 0.288 ;
        RECT 1.8775 0.27 1.8955 0.288 ;
        RECT 1.9855 0.27 2.0035 0.288 ;
        RECT 2.0935 0.27 2.1115 0.288 ;
        RECT 2.284 0.27 2.302 0.288 ;
        RECT 2.353 0.27 2.371 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.53 0.13 1.548 0.159 ;
        RECT 0.882 0.189 1.113 0.207 ;
        RECT 0.882 0.135 0.9 0.207 ;
        RECT 0.558 0.135 0.576 0.165 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 1.093 0.189 1.548 0.207 ;
        RECT 1.53 0.133 1.548 0.207 ;
        RECT 0.882 0.088 0.9 0.155 ;
        RECT 0.558 0.088 0.9 0.106 ;
        RECT 0.234 0.184 0.576 0.202 ;
        RECT 0.558 0.088 0.576 0.202 ;
        RECT 0.234 0.125 0.252 0.202 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
        RECT 0.558 0.137 0.576 0.155 ;
        RECT 0.882 0.137 0.9 0.155 ;
        RECT 1.093 0.189 1.111 0.207 ;
        RECT 1.53 0.133 1.548 0.151 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.682 0.135 1.71 0.153 ;
        RECT 1.044 0.13 1.062 0.16 ;
        RECT 0.72 0.135 0.738 0.165 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 1.6105 0.135 1.708 0.153 ;
        RECT 0.072 0.225 1.6285 0.243 ;
        RECT 1.6105 0.135 1.6285 0.243 ;
        RECT 1.044 0.137 1.062 0.243 ;
        RECT 0.72 0.137 0.738 0.243 ;
        RECT 0.072 0.125 0.09 0.243 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.72 0.137 0.738 0.155 ;
        RECT 1.044 0.137 1.062 0.155 ;
        RECT 1.69 0.135 1.708 0.153 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.854 0.123 1.872 0.153 ;
        RECT 1.206 0.126 1.224 0.158 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 1.854 0.052 1.872 0.151 ;
        RECT 0.396 0.052 1.872 0.07 ;
        RECT 1.206 0.052 1.224 0.151 ;
        RECT 0.396 0.052 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
        RECT 1.206 0.133 1.224 0.151 ;
        RECT 1.854 0.133 1.872 0.151 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.043 0.234 2.196 0.252 ;
        RECT 2.178 0.036 2.196 0.252 ;
        RECT 2.043 0.036 2.196 0.054 ;
      LAYER M2 ;
        RECT 2.178 0.125 2.196 0.158 ;
      LAYER M3 ;
        RECT 2.178 0.126 2.196 0.158 ;
      LAYER V1 ;
        RECT 2.178 0.13 2.196 0.148 ;
      LAYER V2 ;
        RECT 2.178 0.135 2.196 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 1.395 0.1875 1.6735 0.2055 ;
      RECT 1.422 0.0825 1.44 0.2055 ;
      RECT 1.395 0.0825 1.629 0.1005 ;
      RECT 0.018 0.19 0.657 0.208 ;
      RECT 0.018 0.0815 0.036 0.208 ;
      RECT 1.314 0.135 1.386 0.153 ;
      RECT 1.314 0.0815 1.332 0.153 ;
      RECT 0.018 0.0815 1.332 0.0995 ;
      RECT 2.016 0.135 2.034 0.165 ;
      RECT 1.719 0.0795 1.953 0.0975 ;
      RECT 1.719 0.1875 1.953 0.2055 ;
      RECT 1.557 0.0405 1.791 0.0585 ;
      RECT 1.557 0.2295 1.791 0.2475 ;
      RECT 0.909 0.0405 1.467 0.0585 ;
      RECT 0.909 0.2295 1.467 0.2475 ;
      RECT 0.585 0.0405 0.819 0.0585 ;
      RECT 0.585 0.2295 0.819 0.2475 ;
      RECT 0.045 0.0405 0.495 0.0585 ;
      RECT 0.045 0.2295 0.495 0.2475 ;
    LAYER M2 ;
      RECT 1.6535 0.1875 2.034 0.2055 ;
      RECT 2.016 0.137 2.034 0.2055 ;
    LAYER V1 ;
      RECT 2.016 0.137 2.034 0.155 ;
      RECT 1.6535 0.1875 1.6715 0.2055 ;
  END
END MS_3x

MACRO MS_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MS_5x 0 0 ;
  SIZE 3.78 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 3.78 0.018 ;
      LAYER M2 ;
        RECT 0 0 3.78 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.909 0 0.927 0.018 ;
        RECT 1.428 0 1.446 0.018 ;
        RECT 1.9625 0 1.9805 0.018 ;
        RECT 2.259 0 2.277 0.018 ;
        RECT 2.529 0 2.547 0.018 ;
        RECT 2.77 0 2.788 0.018 ;
        RECT 3.339 0 3.357 0.018 ;
        RECT 3.447 0 3.465 0.018 ;
        RECT 3.688 0 3.706 0.018 ;
        RECT 3.757 0 3.775 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 3.78 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 3.78 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.9055 0.27 0.9235 0.288 ;
        RECT 1.1755 0.27 1.1935 0.288 ;
        RECT 1.2835 0.27 1.3015 0.288 ;
        RECT 1.3915 0.27 1.4095 0.288 ;
        RECT 1.4995 0.27 1.5175 0.288 ;
        RECT 1.6075 0.27 1.6255 0.288 ;
        RECT 1.7155 0.27 1.7335 0.288 ;
        RECT 1.8235 0.27 1.8415 0.288 ;
        RECT 1.9315 0.27 1.9495 0.288 ;
        RECT 2.0395 0.27 2.0575 0.288 ;
        RECT 2.0935 0.27 2.1115 0.288 ;
        RECT 2.1475 0.27 2.1655 0.288 ;
        RECT 2.2015 0.27 2.2195 0.288 ;
        RECT 2.3095 0.27 2.3275 0.288 ;
        RECT 2.4175 0.27 2.4355 0.288 ;
        RECT 2.5255 0.27 2.5435 0.288 ;
        RECT 2.77 0.27 2.788 0.288 ;
        RECT 3.0655 0.27 3.0835 0.288 ;
        RECT 3.1735 0.27 3.1915 0.288 ;
        RECT 3.2815 0.27 3.2995 0.288 ;
        RECT 3.3895 0.27 3.4075 0.288 ;
        RECT 3.4975 0.27 3.5155 0.288 ;
        RECT 3.688 0.27 3.706 0.288 ;
        RECT 3.757 0.27 3.775 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.502 0.13 2.52 0.159 ;
        RECT 1.422 0.189 1.761 0.207 ;
        RECT 1.422 0.135 1.44 0.207 ;
        RECT 0.882 0.135 0.9 0.165 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 1.741 0.189 2.52 0.207 ;
        RECT 2.502 0.133 2.52 0.207 ;
        RECT 1.422 0.088 1.44 0.155 ;
        RECT 0.882 0.088 1.44 0.106 ;
        RECT 0.342 0.184 0.9 0.202 ;
        RECT 0.882 0.088 0.9 0.202 ;
        RECT 0.342 0.125 0.36 0.202 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
        RECT 0.882 0.137 0.9 0.155 ;
        RECT 1.422 0.137 1.44 0.155 ;
        RECT 1.741 0.189 1.759 0.207 ;
        RECT 2.502 0.133 2.52 0.151 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.654 0.135 2.79 0.153 ;
        RECT 1.692 0.13 1.71 0.16 ;
        RECT 1.152 0.135 1.17 0.165 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 2.5825 0.135 2.788 0.153 ;
        RECT 0.072 0.225 2.6005 0.243 ;
        RECT 2.5825 0.135 2.6005 0.243 ;
        RECT 1.692 0.137 1.71 0.243 ;
        RECT 1.152 0.137 1.17 0.243 ;
        RECT 0.072 0.125 0.09 0.243 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 1.152 0.137 1.17 0.155 ;
        RECT 1.692 0.137 1.71 0.155 ;
        RECT 2.77 0.135 2.788 0.153 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.042 0.123 3.06 0.153 ;
        RECT 1.962 0.126 1.98 0.158 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 3.042 0.052 3.06 0.151 ;
        RECT 0.612 0.052 3.06 0.07 ;
        RECT 1.962 0.052 1.98 0.151 ;
        RECT 0.612 0.052 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
        RECT 1.962 0.133 1.98 0.151 ;
        RECT 3.042 0.133 3.06 0.151 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.339 0.234 3.6 0.252 ;
        RECT 3.582 0.036 3.6 0.252 ;
        RECT 3.339 0.036 3.6 0.054 ;
      LAYER M2 ;
        RECT 3.582 0.125 3.6 0.158 ;
      LAYER M3 ;
        RECT 3.582 0.126 3.6 0.158 ;
      LAYER V1 ;
        RECT 3.582 0.13 3.6 0.148 ;
      LAYER V2 ;
        RECT 3.582 0.135 3.6 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 2.259 0.1875 2.7555 0.2055 ;
      RECT 2.286 0.0825 2.304 0.2055 ;
      RECT 2.259 0.0825 2.709 0.1005 ;
      RECT 0.018 0.19 1.089 0.208 ;
      RECT 0.018 0.0815 0.036 0.208 ;
      RECT 2.07 0.135 2.25 0.153 ;
      RECT 2.07 0.0815 2.088 0.153 ;
      RECT 0.018 0.0815 2.088 0.0995 ;
      RECT 3.312 0.135 3.33 0.165 ;
      RECT 2.799 0.0795 3.249 0.0975 ;
      RECT 2.799 0.1875 3.249 0.2055 ;
      RECT 2.529 0.0405 2.979 0.0585 ;
      RECT 2.529 0.2295 2.979 0.2475 ;
      RECT 1.449 0.0405 2.439 0.0585 ;
      RECT 1.449 0.2295 2.439 0.2475 ;
      RECT 0.909 0.0405 1.359 0.0585 ;
      RECT 0.909 0.2295 1.359 0.2475 ;
      RECT 0.045 0.0405 0.819 0.0585 ;
      RECT 0.045 0.2295 0.819 0.2475 ;
    LAYER M2 ;
      RECT 2.7355 0.1875 3.33 0.2055 ;
      RECT 3.312 0.137 3.33 0.2055 ;
    LAYER V1 ;
      RECT 3.312 0.137 3.33 0.155 ;
      RECT 2.7355 0.1875 2.7535 0.2055 ;
  END
END MS_5x

MACRO MUX_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX_1x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.348 0 0.366 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
        RECT 0.4505 0 0.4685 0.018 ;
        RECT 0.51 0 0.528 0.018 ;
        RECT 0.546 0 0.564 0.018 ;
        RECT 0.5825 0 0.6005 0.018 ;
        RECT 0.6185 0 0.6365 0.018 ;
        RECT 0.6665 0 0.6845 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.3415 0.27 0.3595 0.288 ;
        RECT 0.393 0.27 0.411 0.288 ;
        RECT 0.44 0.27 0.458 0.288 ;
        RECT 0.51 0.27 0.528 0.288 ;
        RECT 0.546 0.27 0.564 0.288 ;
        RECT 0.5825 0.27 0.6005 0.288 ;
        RECT 0.6185 0.27 0.6365 0.288 ;
        RECT 0.6665 0.27 0.6845 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.585 0.232 0.63 0.25 ;
        RECT 0.612 0.037 0.63 0.25 ;
        RECT 0.585 0.037 0.63 0.055 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END OUT
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.134 0.414 0.164 ;
        RECT 0.288 0.1335 0.306 0.164 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.184 0.414 0.202 ;
        RECT 0.396 0.141 0.414 0.202 ;
        RECT 0.288 0.142 0.306 0.202 ;
        RECT 0.072 0.125 0.09 0.202 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.288 0.142 0.306 0.16 ;
        RECT 0.396 0.141 0.414 0.159 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 0.369 0.232 0.495 0.25 ;
      RECT 0.451 0.037 0.469 0.25 ;
      RECT 0.423 0.037 0.495 0.055 ;
      RECT 0.234 0.189 0.333 0.207 ;
      RECT 0.234 0.08 0.252 0.207 ;
      RECT 0.234 0.08 0.424 0.098 ;
      RECT 0.153 0.232 0.279 0.25 ;
      RECT 0.18 0.037 0.198 0.25 ;
      RECT 0.153 0.037 0.333 0.055 ;
      RECT 0.018 0.232 0.063 0.25 ;
      RECT 0.018 0.056 0.036 0.25 ;
      RECT 0.018 0.056 0.063 0.074 ;
      RECT 0.558 0.078 0.576 0.153 ;
      RECT 0.342 0.123 0.36 0.153 ;
    LAYER M2 ;
      RECT 0.342 0.056 0.36 0.146 ;
      RECT 0.043 0.056 0.36 0.074 ;
      RECT 0.404 0.08 0.576 0.098 ;
    LAYER V1 ;
      RECT 0.558 0.08 0.576 0.098 ;
      RECT 0.404 0.08 0.422 0.098 ;
      RECT 0.342 0.128 0.36 0.146 ;
      RECT 0.043 0.056 0.061 0.074 ;
  END
END MUX_1x

MACRO MUX_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX_2x 0 0 ;
  SIZE 1.188 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.188 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.188 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.061 0 0.079 0.018 ;
        RECT 0.169 0 0.187 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.295 0 0.313 0.018 ;
        RECT 0.3325 0 0.3505 0.018 ;
        RECT 0.369 0 0.387 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
        RECT 0.6665 0 0.6845 0.018 ;
        RECT 0.924 0 0.942 0.018 ;
        RECT 0.984 0 1.002 0.018 ;
        RECT 1.0505 0 1.0685 0.018 ;
        RECT 1.0985 0 1.1165 0.018 ;
        RECT 1.165 0 1.183 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.188 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.188 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.059 0.27 0.077 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.293 0.27 0.311 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.3655 0.27 0.3835 0.288 ;
        RECT 0.5035 0.27 0.5215 0.288 ;
        RECT 0.609 0.27 0.627 0.288 ;
        RECT 0.656 0.27 0.674 0.288 ;
        RECT 0.816 0.27 0.834 0.288 ;
        RECT 1.0145 0.27 1.0325 0.288 ;
        RECT 1.0505 0.27 1.0685 0.288 ;
        RECT 1.0985 0.27 1.1165 0.288 ;
        RECT 1.165 0.27 1.183 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.963 0.232 1.062 0.25 ;
        RECT 1.044 0.037 1.062 0.25 ;
        RECT 0.963 0.037 1.062 0.055 ;
      LAYER M2 ;
        RECT 1.044 0.125 1.062 0.158 ;
      LAYER M3 ;
        RECT 1.044 0.126 1.062 0.158 ;
      LAYER V1 ;
        RECT 1.044 0.13 1.062 0.148 ;
      LAYER V2 ;
        RECT 1.044 0.135 1.062 0.153 ;
    END
  END OUT
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.134 0.63 0.164 ;
        RECT 0.396 0.1335 0.414 0.164 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.184 0.63 0.202 ;
        RECT 0.612 0.141 0.63 0.202 ;
        RECT 0.396 0.142 0.414 0.202 ;
        RECT 0.072 0.125 0.09 0.202 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.396 0.142 0.414 0.16 ;
        RECT 0.612 0.141 0.63 0.159 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 0.531 0.232 0.873 0.25 ;
      RECT 0.774 0.037 0.792 0.25 ;
      RECT 0.639 0.037 0.873 0.055 ;
      RECT 0.342 0.189 0.603 0.207 ;
      RECT 0.342 0.08 0.36 0.207 ;
      RECT 0.342 0.08 0.747 0.098 ;
      RECT 0.207 0.232 0.441 0.25 ;
      RECT 0.288 0.037 0.306 0.25 ;
      RECT 0.207 0.037 0.549 0.055 ;
      RECT 0.018 0.232 0.117 0.25 ;
      RECT 0.018 0.056 0.036 0.25 ;
      RECT 0.018 0.056 0.117 0.074 ;
      RECT 0.936 0.125 0.954 0.153 ;
      RECT 0.504 0.123 0.522 0.153 ;
    LAYER M2 ;
      RECT 0.936 0.08 0.954 0.151 ;
      RECT 0.727 0.08 0.954 0.098 ;
      RECT 0.504 0.056 0.522 0.146 ;
      RECT 0.097 0.056 0.522 0.074 ;
    LAYER V1 ;
      RECT 0.936 0.133 0.954 0.151 ;
      RECT 0.727 0.08 0.745 0.098 ;
      RECT 0.504 0.128 0.522 0.146 ;
      RECT 0.097 0.056 0.115 0.074 ;
  END
END MUX_2x

MACRO MUX_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX_3x 0 0 ;
  SIZE 1.512 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.512 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.512 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.4405 0 0.4585 0.018 ;
        RECT 0.477 0 0.495 0.018 ;
        RECT 0.8065 0 0.8245 0.018 ;
        RECT 0.9905 0 1.0085 0.018 ;
        RECT 1.194 0 1.212 0.018 ;
        RECT 1.3745 0 1.3925 0.018 ;
        RECT 1.4225 0 1.4405 0.018 ;
        RECT 1.489 0 1.507 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.512 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.512 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.4735 0.27 0.4915 0.288 ;
        RECT 0.6655 0.27 0.6835 0.288 ;
        RECT 0.825 0.27 0.843 0.288 ;
        RECT 0.98 0.27 0.998 0.288 ;
        RECT 1.194 0.27 1.212 0.288 ;
        RECT 1.3745 0.27 1.3925 0.288 ;
        RECT 1.4225 0.27 1.4405 0.288 ;
        RECT 1.489 0.27 1.507 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.128 1.062 0.158 ;
      LAYER M2 ;
        RECT 1.044 0.125 1.062 0.158 ;
      LAYER M3 ;
        RECT 1.044 0.126 1.062 0.158 ;
      LAYER V1 ;
        RECT 1.044 0.13 1.062 0.148 ;
      LAYER V2 ;
        RECT 1.044 0.135 1.062 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.233 0.232 1.386 0.25 ;
        RECT 1.368 0.037 1.386 0.25 ;
        RECT 1.233 0.037 1.386 0.055 ;
      LAYER M2 ;
        RECT 1.368 0.125 1.386 0.158 ;
      LAYER M3 ;
        RECT 1.368 0.126 1.386 0.158 ;
      LAYER V1 ;
        RECT 1.368 0.13 1.386 0.148 ;
      LAYER V2 ;
        RECT 1.368 0.135 1.386 0.153 ;
    END
  END OUT
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.134 0.846 0.164 ;
        RECT 0.504 0.1335 0.522 0.164 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.184 0.846 0.202 ;
        RECT 0.828 0.141 0.846 0.202 ;
        RECT 0.504 0.142 0.522 0.202 ;
        RECT 0.072 0.125 0.09 0.202 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.504 0.142 0.522 0.16 ;
        RECT 0.828 0.141 0.846 0.159 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 0.693 0.232 1.143 0.25 ;
      RECT 0.991 0.037 1.009 0.25 ;
      RECT 0.855 0.037 1.143 0.055 ;
      RECT 0.45 0.189 0.765 0.207 ;
      RECT 0.45 0.08 0.468 0.207 ;
      RECT 0.45 0.08 0.964 0.098 ;
      RECT 0.261 0.232 0.603 0.25 ;
      RECT 0.396 0.037 0.414 0.25 ;
      RECT 0.261 0.037 0.765 0.055 ;
      RECT 0.018 0.232 0.171 0.25 ;
      RECT 0.018 0.056 0.036 0.25 ;
      RECT 0.018 0.056 0.227 0.074 ;
      RECT 1.206 0.078 1.224 0.153 ;
      RECT 0.666 0.123 0.684 0.153 ;
    LAYER M2 ;
      RECT 0.666 0.056 0.684 0.146 ;
      RECT 0.207 0.056 0.684 0.074 ;
      RECT 0.944 0.08 1.224 0.098 ;
    LAYER V1 ;
      RECT 1.206 0.08 1.224 0.098 ;
      RECT 0.944 0.08 0.962 0.098 ;
      RECT 0.666 0.128 0.684 0.146 ;
      RECT 0.207 0.056 0.225 0.074 ;
  END
END MUX_3x

MACRO MUX_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX_5x 0 0 ;
  SIZE 2.268 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 2.268 0.018 ;
      LAYER M2 ;
        RECT 0 0 2.268 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.619 0 0.637 0.018 ;
        RECT 0.6565 0 0.6745 0.018 ;
        RECT 0.693 0 0.711 0.018 ;
        RECT 1.2385 0 1.2565 0.018 ;
        RECT 1.5305 0 1.5485 0.018 ;
        RECT 1.842 0 1.86 0.018 ;
        RECT 2.1305 0 2.1485 0.018 ;
        RECT 2.1785 0 2.1965 0.018 ;
        RECT 2.245 0 2.263 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 2.268 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 2.268 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.617 0.27 0.635 0.288 ;
        RECT 0.653 0.27 0.671 0.288 ;
        RECT 0.6895 0.27 0.7075 0.288 ;
        RECT 0.9895 0.27 1.0075 0.288 ;
        RECT 1.257 0.27 1.275 0.288 ;
        RECT 1.5325 0.27 1.5505 0.288 ;
        RECT 1.842 0.27 1.86 0.288 ;
        RECT 2.1305 0.27 2.1485 0.288 ;
        RECT 2.1785 0.27 2.1965 0.288 ;
        RECT 2.245 0.27 2.263 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.128 1.602 0.158 ;
      LAYER M2 ;
        RECT 1.584 0.125 1.602 0.158 ;
      LAYER M3 ;
        RECT 1.584 0.126 1.602 0.158 ;
      LAYER V1 ;
        RECT 1.584 0.13 1.602 0.148 ;
      LAYER V2 ;
        RECT 1.584 0.135 1.602 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.881 0.232 2.142 0.25 ;
        RECT 2.124 0.037 2.142 0.25 ;
        RECT 1.881 0.037 2.142 0.055 ;
      LAYER M2 ;
        RECT 2.124 0.125 2.142 0.158 ;
      LAYER M3 ;
        RECT 2.124 0.126 2.142 0.158 ;
      LAYER V1 ;
        RECT 2.124 0.13 2.142 0.148 ;
      LAYER V2 ;
        RECT 2.124 0.135 2.142 0.153 ;
    END
  END OUT
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.134 1.278 0.164 ;
        RECT 0.72 0.1335 0.738 0.164 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.184 1.278 0.202 ;
        RECT 1.26 0.141 1.278 0.202 ;
        RECT 0.72 0.142 0.738 0.202 ;
        RECT 0.072 0.125 0.09 0.202 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
        RECT 0.72 0.142 0.738 0.16 ;
        RECT 1.26 0.141 1.278 0.159 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1.017 0.232 1.791 0.25 ;
      RECT 1.531 0.037 1.549 0.25 ;
      RECT 1.287 0.037 1.791 0.055 ;
      RECT 0.666 0.189 1.197 0.207 ;
      RECT 0.666 0.08 0.684 0.207 ;
      RECT 0.666 0.08 1.504 0.098 ;
      RECT 0.369 0.232 0.927 0.25 ;
      RECT 0.612 0.037 0.63 0.25 ;
      RECT 0.369 0.037 1.197 0.055 ;
      RECT 0.018 0.232 0.279 0.25 ;
      RECT 0.018 0.056 0.036 0.25 ;
      RECT 0.018 0.056 0.335 0.074 ;
      RECT 1.854 0.078 1.872 0.153 ;
      RECT 0.99 0.123 1.008 0.153 ;
    LAYER M2 ;
      RECT 0.99 0.056 1.008 0.146 ;
      RECT 0.315 0.056 1.008 0.074 ;
      RECT 1.484 0.08 1.872 0.098 ;
    LAYER V1 ;
      RECT 1.854 0.08 1.872 0.098 ;
      RECT 1.484 0.08 1.502 0.098 ;
      RECT 0.99 0.128 1.008 0.146 ;
      RECT 0.315 0.056 0.333 0.074 ;
  END
END MUX_5x

MACRO NAND2_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_1x 0 0 ;
  SIZE 0.324 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.324 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.324 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.301 0 0.319 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.301 0.27 0.319 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.117 0.247 ;
        RECT 0.018 0.041 0.063 0.059 ;
        RECT 0.018 0.041 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
END NAND2_1x

MACRO NAND2_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_2x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.295 0 0.313 0.018 ;
        RECT 0.3325 0 0.3505 0.018 ;
        RECT 0.369 0 0.387 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.293 0.27 0.311 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.3655 0.27 0.3835 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.279 0.247 ;
        RECT 0.018 0.076 0.117 0.094 ;
        RECT 0.018 0.076 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.04 0.279 0.058 ;
  END
END NAND2_2x

MACRO NAND2_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_3x 0 0 ;
  SIZE 0.54 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.54 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.54 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.4405 0 0.4585 0.018 ;
        RECT 0.477 0 0.495 0.018 ;
        RECT 0.517 0 0.535 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.4735 0.27 0.4915 0.288 ;
        RECT 0.517 0.27 0.535 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.333 0.247 ;
        RECT 0.018 0.076 0.171 0.094 ;
        RECT 0.018 0.076 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.099 0.04 0.333 0.058 ;
  END
END NAND2_3x

MACRO NAND2_4x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_4x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.313 0 0.331 0.018 ;
        RECT 0.421 0 0.439 0.018 ;
        RECT 0.511 0 0.529 0.018 ;
        RECT 0.5485 0 0.5665 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.509 0.27 0.527 0.288 ;
        RECT 0.545 0.27 0.563 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.128 0.306 0.158 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.495 0.247 ;
        RECT 0.018 0.076 0.225 0.094 ;
        RECT 0.018 0.076 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.04 0.495 0.058 ;
  END
END NAND2_4x

MACRO NAND2_6x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_6x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.421 0 0.439 0.018 ;
        RECT 0.529 0 0.547 0.018 ;
        RECT 0.637 0 0.655 0.018 ;
        RECT 0.727 0 0.745 0.018 ;
        RECT 0.7645 0 0.7825 0.018 ;
        RECT 0.801 0 0.819 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.527 0.27 0.545 0.288 ;
        RECT 0.635 0.27 0.653 0.288 ;
        RECT 0.725 0.27 0.743 0.288 ;
        RECT 0.761 0.27 0.779 0.288 ;
        RECT 0.7975 0.27 0.8155 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.711 0.247 ;
        RECT 0.018 0.076 0.333 0.094 ;
        RECT 0.018 0.076 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.04 0.711 0.058 ;
  END
END NAND2_6x

MACRO NAND2_8x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_8x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.529 0 0.547 0.018 ;
        RECT 0.637 0 0.655 0.018 ;
        RECT 0.745 0 0.763 0.018 ;
        RECT 0.853 0 0.871 0.018 ;
        RECT 0.943 0 0.961 0.018 ;
        RECT 0.9805 0 0.9985 0.018 ;
        RECT 1.017 0 1.035 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.527 0.27 0.545 0.288 ;
        RECT 0.635 0.27 0.653 0.288 ;
        RECT 0.743 0.27 0.761 0.288 ;
        RECT 0.851 0.27 0.869 0.288 ;
        RECT 0.941 0.27 0.959 0.288 ;
        RECT 0.977 0.27 0.995 0.288 ;
        RECT 1.0135 0.27 1.0315 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.927 0.247 ;
        RECT 0.018 0.076 0.441 0.094 ;
        RECT 0.018 0.076 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.04 0.927 0.058 ;
  END
END NAND2_8x

MACRO NAND3_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_1x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.315 0 0.333 0.018 ;
        RECT 0.351 0 0.369 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.3115 0.27 0.3295 0.288 ;
        RECT 0.3475 0.27 0.3655 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.171 0.247 ;
        RECT 0.018 0.04 0.063 0.058 ;
        RECT 0.018 0.04 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
END NAND3_1x

MACRO NAND3_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_2x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.169 0 0.187 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.531 0 0.549 0.018 ;
        RECT 0.567 0 0.585 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.5275 0.27 0.5455 0.288 ;
        RECT 0.5635 0.27 0.5815 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.441 0.247 ;
        RECT 0.018 0.085 0.117 0.103 ;
        RECT 0.018 0.085 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.207 0.085 0.441 0.103 ;
      RECT 0.045 0.049 0.279 0.067 ;
  END
END NAND3_2x

MACRO NAND3_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_3x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.223 0 0.241 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.639 0 0.657 0.018 ;
        RECT 0.675 0 0.693 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.6355 0.27 0.6535 0.288 ;
        RECT 0.6715 0.27 0.6895 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.495 0.247 ;
        RECT 0.018 0.085 0.171 0.103 ;
        RECT 0.018 0.085 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.261 0.085 0.495 0.103 ;
      RECT 0.099 0.049 0.333 0.067 ;
  END
END NAND3_3x

MACRO NAND3_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_5x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.331 0 0.349 0.018 ;
        RECT 0.619 0 0.637 0.018 ;
        RECT 0.999 0 1.017 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.653 0.27 0.671 0.288 ;
        RECT 0.761 0.27 0.779 0.288 ;
        RECT 0.9955 0.27 1.0135 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.819 0.247 ;
        RECT 0.018 0.085 0.279 0.103 ;
        RECT 0.018 0.085 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.369 0.085 0.819 0.103 ;
      RECT 0.099 0.049 0.549 0.067 ;
  END
END NAND3_5x

MACRO NAND3_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_7x 0 0 ;
  SIZE 1.404 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.404 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.404 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.439 0 0.457 0.018 ;
        RECT 0.835 0 0.853 0.018 ;
        RECT 1.323 0 1.341 0.018 ;
        RECT 1.381 0 1.399 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.404 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.404 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.311 0.27 0.329 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.869 0.27 0.887 0.288 ;
        RECT 0.977 0.27 0.995 0.288 ;
        RECT 1.085 0.27 1.103 0.288 ;
        RECT 1.3195 0.27 1.3375 0.288 ;
        RECT 1.381 0.27 1.399 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 1.143 0.247 ;
        RECT 0.018 0.085 0.387 0.103 ;
        RECT 0.018 0.085 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.477 0.085 1.143 0.103 ;
      RECT 0.099 0.049 0.765 0.067 ;
  END
END NAND3_7x

MACRO NOR2_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_1x 0 0 ;
  SIZE 0.324 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.324 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.324 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.301 0 0.319 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.324 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.301 0.27 0.319 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.153 0.229 0.198 0.247 ;
        RECT 0.18 0.041 0.198 0.247 ;
        RECT 0.099 0.041 0.198 0.059 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END OUT
END NOR2_1x

MACRO NOR2_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_2x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0955 0 0.1135 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.295 0 0.313 0.018 ;
        RECT 0.3325 0 0.3505 0.018 ;
        RECT 0.369 0 0.387 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.068 0.27 0.086 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.293 0.27 0.311 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.3655 0.27 0.3835 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.193 0.306 0.211 ;
        RECT 0.288 0.041 0.306 0.211 ;
        RECT 0.045 0.041 0.306 0.059 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.279 0.247 ;
  END
END NOR2_2x

MACRO NOR2_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_3x 0 0 ;
  SIZE 0.54 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.54 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.54 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.4405 0 0.4585 0.018 ;
        RECT 0.477 0 0.495 0.018 ;
        RECT 0.517 0 0.535 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.068 0.27 0.086 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.401 0.27 0.419 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 0.4735 0.27 0.4915 0.288 ;
        RECT 0.517 0.27 0.535 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.193 0.414 0.211 ;
        RECT 0.396 0.041 0.414 0.211 ;
        RECT 0.099 0.041 0.414 0.059 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.099 0.229 0.333 0.247 ;
  END
END NOR2_3x

MACRO NOR2_4x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_4x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0955 0 0.1135 0.018 ;
        RECT 0.2035 0 0.2215 0.018 ;
        RECT 0.313 0 0.331 0.018 ;
        RECT 0.421 0 0.439 0.018 ;
        RECT 0.511 0 0.529 0.018 ;
        RECT 0.5485 0 0.5665 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.068 0.27 0.086 0.288 ;
        RECT 0.176 0.27 0.194 0.288 ;
        RECT 0.275 0.27 0.293 0.288 ;
        RECT 0.383 0.27 0.401 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.509 0.27 0.527 0.288 ;
        RECT 0.545 0.27 0.563 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.128 0.306 0.158 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.315 0.193 0.522 0.211 ;
        RECT 0.504 0.041 0.522 0.211 ;
        RECT 0.045 0.041 0.522 0.059 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.495 0.247 ;
  END
END NOR2_4x

MACRO NOR2_6x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_6x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0955 0 0.1135 0.018 ;
        RECT 0.2035 0 0.2215 0.018 ;
        RECT 0.3115 0 0.3295 0.018 ;
        RECT 0.421 0 0.439 0.018 ;
        RECT 0.529 0 0.547 0.018 ;
        RECT 0.637 0 0.655 0.018 ;
        RECT 0.727 0 0.745 0.018 ;
        RECT 0.7645 0 0.7825 0.018 ;
        RECT 0.801 0 0.819 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.068 0.27 0.086 0.288 ;
        RECT 0.176 0.27 0.194 0.288 ;
        RECT 0.284 0.27 0.302 0.288 ;
        RECT 0.383 0.27 0.401 0.288 ;
        RECT 0.491 0.27 0.509 0.288 ;
        RECT 0.599 0.27 0.617 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.725 0.27 0.743 0.288 ;
        RECT 0.761 0.27 0.779 0.288 ;
        RECT 0.7975 0.27 0.8155 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.193 0.738 0.211 ;
        RECT 0.72 0.041 0.738 0.211 ;
        RECT 0.045 0.041 0.738 0.059 ;
      LAYER M2 ;
        RECT 0.72 0.125 0.738 0.158 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.711 0.247 ;
  END
END NOR2_6x

MACRO NOR2_8x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_8x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0955 0 0.1135 0.018 ;
        RECT 0.2035 0 0.2215 0.018 ;
        RECT 0.3115 0 0.3295 0.018 ;
        RECT 0.4195 0 0.4375 0.018 ;
        RECT 0.529 0 0.547 0.018 ;
        RECT 0.637 0 0.655 0.018 ;
        RECT 0.745 0 0.763 0.018 ;
        RECT 0.853 0 0.871 0.018 ;
        RECT 0.9805 0 0.9985 0.018 ;
        RECT 1.017 0 1.035 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.068 0.27 0.086 0.288 ;
        RECT 0.176 0.27 0.194 0.288 ;
        RECT 0.284 0.27 0.302 0.288 ;
        RECT 0.3585 0.27 0.3765 0.288 ;
        RECT 0.4665 0.27 0.4845 0.288 ;
        RECT 0.599 0.27 0.617 0.288 ;
        RECT 0.707 0.27 0.725 0.288 ;
        RECT 0.815 0.27 0.833 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 0.977 0.27 0.995 0.288 ;
        RECT 1.0135 0.27 1.0315 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.531 0.193 0.954 0.211 ;
        RECT 0.936 0.041 0.954 0.211 ;
        RECT 0.045 0.041 0.954 0.059 ;
      LAYER M2 ;
        RECT 0.936 0.125 0.954 0.158 ;
      LAYER M3 ;
        RECT 0.936 0.126 0.954 0.158 ;
      LAYER V1 ;
        RECT 0.936 0.13 0.954 0.148 ;
      LAYER V2 ;
        RECT 0.936 0.135 0.954 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.927 0.247 ;
  END
END NOR2_8x

MACRO NOR3_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_1x 0 0 ;
  SIZE 0.378 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.378 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.378 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.241 0 0.259 0.018 ;
        RECT 0.2785 0 0.2965 0.018 ;
        RECT 0.315 0 0.333 0.018 ;
        RECT 0.355 0 0.373 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.378 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.378 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.239 0.27 0.257 0.288 ;
        RECT 0.275 0.27 0.293 0.288 ;
        RECT 0.3115 0.27 0.3295 0.288 ;
        RECT 0.355 0.27 0.373 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.229 0.252 0.247 ;
        RECT 0.234 0.041 0.252 0.247 ;
        RECT 0.099 0.041 0.252 0.059 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END OUT
END NOR3_1x

MACRO NOR3_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_2x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.511 0 0.529 0.018 ;
        RECT 0.5485 0 0.5665 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.095 0.27 0.113 0.288 ;
        RECT 0.167 0.27 0.185 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.509 0.27 0.527 0.288 ;
        RECT 0.545 0.27 0.563 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.185 0.522 0.203 ;
        RECT 0.504 0.041 0.522 0.203 ;
        RECT 0.099 0.041 0.522 0.059 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.207 0.229 0.495 0.247 ;
      RECT 0.045 0.184 0.279 0.202 ;
  END
END NOR3_2x

MACRO NOR3_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_3x 0 0 ;
  SIZE 0.702 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.702 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.702 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.565 0 0.583 0.018 ;
        RECT 0.6025 0 0.6205 0.018 ;
        RECT 0.639 0 0.657 0.018 ;
        RECT 0.679 0 0.697 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.702 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.702 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.527 0.27 0.545 0.288 ;
        RECT 0.563 0.27 0.581 0.288 ;
        RECT 0.599 0.27 0.617 0.288 ;
        RECT 0.6355 0.27 0.6535 0.288 ;
        RECT 0.679 0.27 0.697 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.185 0.576 0.203 ;
        RECT 0.558 0.041 0.576 0.203 ;
        RECT 0.099 0.041 0.576 0.059 ;
      LAYER M2 ;
        RECT 0.558 0.125 0.576 0.158 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.261 0.229 0.495 0.247 ;
      RECT 0.099 0.184 0.333 0.202 ;
  END
END NOR3_3x

MACRO NOR3_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_5x 0 0 ;
  SIZE 1.026 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.026 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.026 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.3655 0 0.3835 0.018 ;
        RECT 0.4735 0 0.4915 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.691 0 0.709 0.018 ;
        RECT 0.799 0 0.817 0.018 ;
        RECT 0.889 0 0.907 0.018 ;
        RECT 0.9265 0 0.9445 0.018 ;
        RECT 0.963 0 0.981 0.018 ;
        RECT 1.003 0 1.021 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.026 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.026 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.329 0.27 0.347 0.288 ;
        RECT 0.851 0.27 0.869 0.288 ;
        RECT 0.887 0.27 0.905 0.288 ;
        RECT 0.923 0.27 0.941 0.288 ;
        RECT 0.9595 0.27 0.9775 0.288 ;
        RECT 1.003 0.27 1.021 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.639 0.185 0.9 0.203 ;
        RECT 0.882 0.041 0.9 0.203 ;
        RECT 0.099 0.041 0.9 0.059 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.369 0.229 0.819 0.247 ;
      RECT 0.099 0.184 0.549 0.202 ;
  END
END NOR3_5x

MACRO NOR3_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_7x 0 0 ;
  SIZE 1.35 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.35 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.35 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.3655 0 0.3835 0.018 ;
        RECT 0.4735 0 0.4915 0.018 ;
        RECT 0.5815 0 0.5995 0.018 ;
        RECT 0.6895 0 0.7075 0.018 ;
        RECT 0.799 0 0.817 0.018 ;
        RECT 0.907 0 0.925 0.018 ;
        RECT 1.015 0 1.033 0.018 ;
        RECT 1.123 0 1.141 0.018 ;
        RECT 1.213 0 1.231 0.018 ;
        RECT 1.2505 0 1.2685 0.018 ;
        RECT 1.287 0 1.305 0.018 ;
        RECT 1.327 0 1.345 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.35 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.35 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.437 0.27 0.455 0.288 ;
        RECT 1.175 0.27 1.193 0.288 ;
        RECT 1.211 0.27 1.229 0.288 ;
        RECT 1.247 0.27 1.265 0.288 ;
        RECT 1.2835 0.27 1.3015 0.288 ;
        RECT 1.327 0.27 1.345 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.185 1.224 0.203 ;
        RECT 1.206 0.041 1.224 0.203 ;
        RECT 0.099 0.041 1.224 0.059 ;
      LAYER M2 ;
        RECT 1.206 0.125 1.224 0.158 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.477 0.229 1.143 0.247 ;
      RECT 0.099 0.184 0.765 0.202 ;
  END
END NOR3_7x


MACRO OAI21_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_1x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.315 0 0.333 0.018 ;
        RECT 0.351 0 0.369 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.3115 0.27 0.3295 0.288 ;
        RECT 0.3475 0.27 0.3655 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.229 0.252 0.247 ;
        RECT 0.234 0.04 0.252 0.247 ;
        RECT 0.207 0.04 0.252 0.058 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 0.171 0.059 ;
  END
END OAI21_1x

MACRO OAI21_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_2x 0 0 ;
  SIZE 0.648 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.648 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.648 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.4945 0 0.5125 0.018 ;
        RECT 0.531 0 0.549 0.018 ;
        RECT 0.567 0 0.585 0.018 ;
        RECT 0.625 0 0.643 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.648 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.491 0.27 0.509 0.288 ;
        RECT 0.5275 0.27 0.5455 0.288 ;
        RECT 0.5635 0.27 0.5815 0.288 ;
        RECT 0.625 0.27 0.643 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.229 0.522 0.247 ;
        RECT 0.504 0.082 0.522 0.247 ;
        RECT 0.423 0.082 0.522 0.1 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 0.495 0.059 ;
      RECT 0.045 0.187 0.279 0.205 ;
  END
END OAI21_2x

MACRO OAI21_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_3x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.5485 0 0.5665 0.018 ;
        RECT 0.639 0 0.657 0.018 ;
        RECT 0.675 0 0.693 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.545 0.27 0.563 0.288 ;
        RECT 0.6715 0.27 0.6895 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.229 0.576 0.247 ;
        RECT 0.558 0.082 0.576 0.247 ;
        RECT 0.423 0.082 0.576 0.1 ;
      LAYER M2 ;
        RECT 0.558 0.125 0.576 0.158 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 0.495 0.059 ;
      RECT 0.099 0.187 0.333 0.205 ;
  END
END OAI21_3x

MACRO OAI21_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_5x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.8725 0 0.8905 0.018 ;
        RECT 0.963 0 0.981 0.018 ;
        RECT 0.999 0 1.017 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.869 0.27 0.887 0.288 ;
        RECT 0.9595 0.27 0.9775 0.288 ;
        RECT 0.9955 0.27 1.0135 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.229 0.9 0.247 ;
        RECT 0.882 0.082 0.9 0.247 ;
        RECT 0.639 0.082 0.9 0.1 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 0.819 0.059 ;
      RECT 0.099 0.187 0.549 0.205 ;
  END
END OAI21_5x

MACRO OAI21_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_7x 0 0 ;
  SIZE 1.404 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.404 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.404 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 1.1965 0 1.2145 0.018 ;
        RECT 1.287 0 1.305 0.018 ;
        RECT 1.323 0 1.341 0.018 ;
        RECT 1.381 0 1.399 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.404 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.404 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.193 0.27 1.211 0.288 ;
        RECT 1.2835 0.27 1.3015 0.288 ;
        RECT 1.3195 0.27 1.3375 0.288 ;
        RECT 1.381 0.27 1.399 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.229 1.224 0.247 ;
        RECT 1.206 0.082 1.224 0.247 ;
        RECT 0.855 0.082 1.224 0.1 ;
      LAYER M2 ;
        RECT 1.206 0.125 1.224 0.158 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 1.143 0.059 ;
      RECT 0.099 0.187 0.765 0.205 ;
  END
END OAI21_7x

MACRO OAI22_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_1x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.348 0 0.366 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.3415 0.27 0.3595 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.229 0.279 0.247 ;
        RECT 0.018 0.082 0.117 0.1 ;
        RECT 0.018 0.082 0.036 0.247 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 0.279 0.059 ;
  END
END OAI22_1x

MACRO OAI22_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_2x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.511 0 0.529 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.621 0 0.639 0.018 ;
        RECT 0.672 0 0.69 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.6175 0.27 0.6355 0.288 ;
        RECT 0.6655 0.27 0.6835 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.183 0.549 0.201 ;
        RECT 0.018 0.082 0.279 0.1 ;
        RECT 0.018 0.082 0.036 0.201 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.369 0.226 0.603 0.244 ;
      RECT 0.099 0.041 0.549 0.059 ;
      RECT 0.045 0.226 0.279 0.244 ;
  END
END OAI22_2x

MACRO OAI22_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_3x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.565 0 0.583 0.018 ;
        RECT 0.639 0 0.657 0.018 ;
        RECT 0.729 0 0.747 0.018 ;
        RECT 0.78 0 0.798 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.6895 0.27 0.7075 0.288 ;
        RECT 0.7255 0.27 0.7435 0.288 ;
        RECT 0.7735 0.27 0.7915 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.128 0.576 0.158 ;
      LAYER M2 ;
        RECT 0.558 0.125 0.576 0.158 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.183 0.711 0.201 ;
        RECT 0.018 0.082 0.333 0.1 ;
        RECT 0.018 0.082 0.036 0.201 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 0.711 0.059 ;
      RECT 0.423 0.226 0.657 0.244 ;
      RECT 0.099 0.226 0.333 0.244 ;
  END
END OAI22_3x

MACRO OAI22_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_5x 0 0 ;
  SIZE 1.296 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.296 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.296 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.619 0 0.637 0.018 ;
        RECT 0.889 0 0.907 0.018 ;
        RECT 0.963 0 0.981 0.018 ;
        RECT 1.071 0 1.089 0.018 ;
        RECT 1.161 0 1.179 0.018 ;
        RECT 1.212 0 1.23 0.018 ;
        RECT 1.273 0 1.291 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 1.1215 0.27 1.1395 0.288 ;
        RECT 1.1575 0.27 1.1755 0.288 ;
        RECT 1.2055 0.27 1.2235 0.288 ;
        RECT 1.273 0.27 1.291 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.882 0.128 0.9 0.158 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.183 1.143 0.201 ;
        RECT 0.018 0.082 0.549 0.1 ;
        RECT 0.018 0.082 0.036 0.201 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 1.143 0.059 ;
      RECT 0.639 0.226 1.089 0.244 ;
      RECT 0.099 0.226 0.549 0.244 ;
  END
END OAI22_5x

MACRO OAI22_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_7x 0 0 ;
  SIZE 1.728 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.728 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.728 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.835 0 0.853 0.018 ;
        RECT 1.213 0 1.231 0.018 ;
        RECT 1.287 0 1.305 0.018 ;
        RECT 1.395 0 1.413 0.018 ;
        RECT 1.503 0 1.521 0.018 ;
        RECT 1.593 0 1.611 0.018 ;
        RECT 1.644 0 1.662 0.018 ;
        RECT 1.705 0 1.723 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.5895 0.27 1.6075 0.288 ;
        RECT 1.6375 0.27 1.6555 0.288 ;
        RECT 1.705 0.27 1.723 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.128 1.224 0.158 ;
      LAYER M2 ;
        RECT 1.206 0.125 1.224 0.158 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.183 1.575 0.201 ;
        RECT 0.018 0.082 0.765 0.1 ;
        RECT 0.018 0.082 0.036 0.201 ;
      LAYER M2 ;
        RECT 0.018 0.125 0.036 0.158 ;
      LAYER M3 ;
        RECT 0.018 0.126 0.036 0.158 ;
      LAYER V1 ;
        RECT 0.018 0.13 0.036 0.148 ;
      LAYER V2 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.041 1.575 0.059 ;
      RECT 0.855 0.226 1.521 0.244 ;
      RECT 0.099 0.226 0.765 0.244 ;
  END
END OAI22_7x

MACRO OAOI211_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211_1x 0 0 ;
  SIZE 0.432 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.432 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.333 0 0.351 0.018 ;
        RECT 0.409 0 0.427 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.432 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.33 0.27 0.348 0.288 ;
        RECT 0.366 0.27 0.384 0.288 ;
        RECT 0.409 0.27 0.427 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.128 0.144 0.158 ;
      LAYER M2 ;
        RECT 0.126 0.125 0.144 0.158 ;
      LAYER M3 ;
        RECT 0.126 0.126 0.144 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.13 0.144 0.148 ;
      LAYER V2 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.189 0.306 0.207 ;
        RECT 0.288 0.085 0.306 0.207 ;
        RECT 0.099 0.085 0.306 0.103 ;
      LAYER M2 ;
        RECT 0.288 0.125 0.306 0.158 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.225 0.247 ;
      RECT 0.045 0.042 0.171 0.06 ;
  END
END OAOI211_1x

MACRO OAOI211_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211_2x 0 0 ;
  SIZE 0.756 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.756 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.756 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.621 0 0.639 0.018 ;
        RECT 0.657 0 0.675 0.018 ;
        RECT 0.733 0 0.751 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.756 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.6175 0.27 0.6355 0.288 ;
        RECT 0.654 0.27 0.672 0.288 ;
        RECT 0.69 0.27 0.708 0.288 ;
        RECT 0.733 0.27 0.751 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.128 0.198 0.158 ;
      LAYER M2 ;
        RECT 0.18 0.125 0.198 0.158 ;
      LAYER M3 ;
        RECT 0.18 0.126 0.198 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.13 0.198 0.148 ;
      LAYER V2 ;
        RECT 0.18 0.135 0.198 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
      LAYER M2 ;
        RECT 0.504 0.125 0.522 0.158 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.531 0.189 0.63 0.207 ;
        RECT 0.612 0.085 0.63 0.207 ;
        RECT 0.045 0.085 0.63 0.103 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.477 0.234 0.603 0.252 ;
      RECT 0.477 0.186 0.495 0.252 ;
      RECT 0.099 0.186 0.495 0.204 ;
      RECT 0.099 0.042 0.441 0.06 ;
      RECT 0.045 0.229 0.279 0.247 ;
  END
END OAOI211_2x

MACRO OAOI211_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211_3x 0 0 ;
  SIZE 0.864 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.864 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.403 0 0.421 0.018 ;
        RECT 0.639 0 0.657 0.018 ;
        RECT 0.729 0 0.747 0.018 ;
        RECT 0.765 0 0.783 0.018 ;
        RECT 0.841 0 0.859 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.864 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.6895 0.27 0.7075 0.288 ;
        RECT 0.7255 0.27 0.7435 0.288 ;
        RECT 0.762 0.27 0.78 0.288 ;
        RECT 0.798 0.27 0.816 0.288 ;
        RECT 0.841 0.27 0.859 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
      LAYER M2 ;
        RECT 0.234 0.125 0.252 0.158 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.128 0.414 0.158 ;
      LAYER M2 ;
        RECT 0.396 0.125 0.414 0.158 ;
      LAYER M3 ;
        RECT 0.396 0.126 0.414 0.158 ;
      LAYER V1 ;
        RECT 0.396 0.13 0.414 0.148 ;
      LAYER V2 ;
        RECT 0.396 0.135 0.414 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.128 0.576 0.158 ;
      LAYER M2 ;
        RECT 0.558 0.125 0.576 0.158 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.585 0.189 0.738 0.207 ;
        RECT 0.72 0.085 0.738 0.207 ;
        RECT 0.099 0.085 0.738 0.103 ;
      LAYER M2 ;
        RECT 0.72 0.125 0.738 0.158 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 0.657 0.247 ;
      RECT 0.045 0.042 0.495 0.06 ;
      RECT 0.099 0.186 0.333 0.204 ;
  END
END OAOI211_3x

MACRO OAOI211_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211_5x 0 0 ;
  SIZE 1.296 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.296 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.296 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.619 0 0.637 0.018 ;
        RECT 0.963 0 0.981 0.018 ;
        RECT 1.071 0 1.089 0.018 ;
        RECT 1.161 0 1.179 0.018 ;
        RECT 1.197 0 1.215 0.018 ;
        RECT 1.273 0 1.291 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.296 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 1.1215 0.27 1.1395 0.288 ;
        RECT 1.1575 0.27 1.1755 0.288 ;
        RECT 1.194 0.27 1.212 0.288 ;
        RECT 1.23 0.27 1.248 0.288 ;
        RECT 1.273 0.27 1.291 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.128 0.36 0.158 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.128 0.63 0.158 ;
      LAYER M2 ;
        RECT 0.612 0.125 0.63 0.158 ;
      LAYER M3 ;
        RECT 0.612 0.126 0.63 0.158 ;
      LAYER V1 ;
        RECT 0.612 0.13 0.63 0.148 ;
      LAYER V2 ;
        RECT 0.612 0.135 0.63 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.882 0.128 0.9 0.158 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.909 0.189 1.17 0.207 ;
        RECT 1.152 0.085 1.17 0.207 ;
        RECT 0.099 0.085 1.17 0.103 ;
      LAYER M2 ;
        RECT 1.152 0.125 1.17 0.158 ;
      LAYER M3 ;
        RECT 1.152 0.126 1.17 0.158 ;
      LAYER V1 ;
        RECT 1.152 0.13 1.17 0.148 ;
      LAYER V2 ;
        RECT 1.152 0.135 1.17 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 1.089 0.247 ;
      RECT 0.045 0.042 0.819 0.06 ;
      RECT 0.099 0.186 0.549 0.204 ;
  END
END OAOI211_5x

MACRO OAOI211_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211_7x 0 0 ;
  SIZE 1.728 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.728 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.728 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.835 0 0.853 0.018 ;
        RECT 1.287 0 1.305 0.018 ;
        RECT 1.395 0 1.413 0.018 ;
        RECT 1.503 0 1.521 0.018 ;
        RECT 1.593 0 1.611 0.018 ;
        RECT 1.629 0 1.647 0.018 ;
        RECT 1.705 0 1.723 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.728 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.5535 0.27 1.5715 0.288 ;
        RECT 1.5895 0.27 1.6075 0.288 ;
        RECT 1.626 0.27 1.644 0.288 ;
        RECT 1.662 0.27 1.68 0.288 ;
        RECT 1.705 0.27 1.723 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.128 0.468 0.158 ;
      LAYER M2 ;
        RECT 0.45 0.125 0.468 0.158 ;
      LAYER M3 ;
        RECT 0.45 0.126 0.468 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.13 0.468 0.148 ;
      LAYER V2 ;
        RECT 0.45 0.135 0.468 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.128 0.09 0.158 ;
      LAYER M2 ;
        RECT 0.072 0.125 0.09 0.158 ;
      LAYER M3 ;
        RECT 0.072 0.126 0.09 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.13 0.09 0.148 ;
      LAYER V2 ;
        RECT 0.072 0.135 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.128 0.846 0.158 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.128 1.224 0.158 ;
      LAYER M2 ;
        RECT 1.206 0.125 1.224 0.158 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.233 0.189 1.602 0.207 ;
        RECT 1.584 0.085 1.602 0.207 ;
        RECT 0.099 0.085 1.602 0.103 ;
      LAYER M2 ;
        RECT 1.584 0.125 1.602 0.158 ;
      LAYER M3 ;
        RECT 1.584 0.126 1.602 0.158 ;
      LAYER V1 ;
        RECT 1.584 0.13 1.602 0.148 ;
      LAYER V2 ;
        RECT 1.584 0.135 1.602 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.045 0.229 1.521 0.247 ;
      RECT 0.045 0.042 1.143 0.06 ;
      RECT 0.099 0.186 0.765 0.204 ;
  END
END OAOI211_7x

MACRO XNOR2_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_1x 0 0 ;
  SIZE 0.54 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.54 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.54 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.115 0 0.133 0.018 ;
        RECT 0.151 0 0.169 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.348 0 0.366 0.018 ;
        RECT 0.4505 0 0.4685 0.018 ;
        RECT 0.517 0 0.535 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.3415 0.27 0.3595 0.288 ;
        RECT 0.4435 0.27 0.4615 0.288 ;
        RECT 0.517 0.27 0.535 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.128 0.306 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 0.306 0.232 ;
        RECT 0.288 0.125 0.306 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
        RECT 0.126 0.132 0.144 0.162 ;
      LAYER M2 ;
        RECT 0.126 0.178 0.252 0.196 ;
        RECT 0.234 0.125 0.252 0.196 ;
        RECT 0.126 0.134 0.144 0.196 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.139 0.144 0.157 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.229 0.36 0.247 ;
        RECT 0.342 0.085 0.36 0.247 ;
        RECT 0.261 0.085 0.36 0.103 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.117 0.247 ;
      RECT 0.018 0.0865 0.036 0.247 ;
      RECT 0.18 0.0865 0.198 0.15 ;
      RECT 0.018 0.0865 0.198 0.1045 ;
      RECT 0.207 0.042 0.333 0.06 ;
  END
END XNOR2_1x

MACRO XNOR2_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_2x 0 0 ;
  SIZE 0.972 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.972 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.972 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.169 0 0.187 0.018 ;
        RECT 0.205 0 0.223 0.018 ;
        RECT 0.421 0 0.439 0.018 ;
        RECT 0.4945 0 0.5125 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.834 0 0.852 0.018 ;
        RECT 0.8825 0 0.9005 0.018 ;
        RECT 0.949 0 0.967 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.972 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.972 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.491 0.27 0.509 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.8275 0.27 0.8455 0.288 ;
        RECT 0.8755 0.27 0.8935 0.288 ;
        RECT 0.949 0.27 0.967 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.128 0.738 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 0.738 0.232 ;
        RECT 0.72 0.125 0.738 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
        RECT 0.18 0.132 0.198 0.162 ;
      LAYER M2 ;
        RECT 0.18 0.178 0.522 0.196 ;
        RECT 0.504 0.125 0.522 0.196 ;
        RECT 0.18 0.134 0.198 0.196 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.139 0.198 0.157 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.369 0.185 0.846 0.203 ;
        RECT 0.828 0.085 0.846 0.203 ;
        RECT 0.531 0.085 0.846 0.103 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.225 0.247 ;
      RECT 0.018 0.0865 0.036 0.247 ;
      RECT 0.396 0.0865 0.414 0.15 ;
      RECT 0.018 0.0865 0.414 0.1045 ;
      RECT 0.531 0.228 0.819 0.246 ;
      RECT 0.369 0.042 0.765 0.06 ;
      RECT 0.045 0.042 0.279 0.06 ;
  END
END XNOR2_2x

MACRO XNOR2_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_3x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.259 0 0.277 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.5485 0 0.5665 0.018 ;
        RECT 0.693 0 0.711 0.018 ;
        RECT 0.888 0 0.906 0.018 ;
        RECT 0.9905 0 1.0085 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.545 0.27 0.563 0.288 ;
        RECT 0.6895 0.27 0.7075 0.288 ;
        RECT 0.8815 0.27 0.8995 0.288 ;
        RECT 0.9835 0.27 1.0015 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.128 0.738 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 0.738 0.232 ;
        RECT 0.72 0.125 0.738 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.128 0.576 0.158 ;
        RECT 0.234 0.132 0.252 0.162 ;
      LAYER M2 ;
        RECT 0.234 0.178 0.576 0.196 ;
        RECT 0.558 0.125 0.576 0.196 ;
        RECT 0.234 0.134 0.252 0.196 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.139 0.252 0.157 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.185 0.9 0.203 ;
        RECT 0.882 0.085 0.9 0.203 ;
        RECT 0.585 0.085 0.9 0.103 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.333 0.247 ;
      RECT 0.018 0.0865 0.036 0.247 ;
      RECT 0.396 0.0865 0.414 0.15 ;
      RECT 0.018 0.0865 0.414 0.1045 ;
      RECT 0.423 0.042 0.873 0.06 ;
      RECT 0.585 0.228 0.819 0.246 ;
      RECT 0.099 0.042 0.333 0.06 ;
  END
END XNOR2_3x

MACRO XNOR2_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_5x 0 0 ;
  SIZE 1.62 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.62 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.62 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.367 0 0.385 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.691 0 0.709 0.018 ;
        RECT 0.799 0 0.817 0.018 ;
        RECT 0.8725 0 0.8905 0.018 ;
        RECT 1.125 0 1.143 0.018 ;
        RECT 1.428 0 1.446 0.018 ;
        RECT 1.5305 0 1.5485 0.018 ;
        RECT 1.597 0 1.615 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.62 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.62 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.869 0.27 0.887 0.288 ;
        RECT 1.1215 0.27 1.1395 0.288 ;
        RECT 1.4215 0.27 1.4395 0.288 ;
        RECT 1.5235 0.27 1.5415 0.288 ;
        RECT 1.597 0.27 1.615 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.128 1.17 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 1.17 0.232 ;
        RECT 1.152 0.125 1.17 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 1.152 0.126 1.17 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 1.152 0.13 1.17 0.148 ;
      LAYER V2 ;
        RECT 1.152 0.135 1.17 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.882 0.128 0.9 0.158 ;
        RECT 0.342 0.132 0.36 0.162 ;
      LAYER M2 ;
        RECT 0.342 0.178 0.9 0.196 ;
        RECT 0.882 0.125 0.9 0.196 ;
        RECT 0.342 0.134 0.36 0.196 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.139 0.36 0.157 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.639 0.185 1.44 0.203 ;
        RECT 1.422 0.085 1.44 0.203 ;
        RECT 0.909 0.085 1.44 0.103 ;
      LAYER M2 ;
        RECT 1.422 0.125 1.44 0.158 ;
      LAYER M3 ;
        RECT 1.422 0.126 1.44 0.158 ;
      LAYER V1 ;
        RECT 1.422 0.13 1.44 0.148 ;
      LAYER V2 ;
        RECT 1.422 0.135 1.44 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.549 0.247 ;
      RECT 0.018 0.0865 0.036 0.247 ;
      RECT 0.612 0.0865 0.63 0.15 ;
      RECT 0.018 0.0865 0.63 0.1045 ;
      RECT 0.639 0.042 1.413 0.06 ;
      RECT 0.909 0.228 1.359 0.246 ;
      RECT 0.099 0.042 0.549 0.06 ;
  END
END XNOR2_5x

MACRO XNOR2_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_7x 0 0 ;
  SIZE 2.16 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 2.16 0.018 ;
      LAYER M2 ;
        RECT 0 0 2.16 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.475 0 0.493 0.018 ;
        RECT 0.583 0 0.601 0.018 ;
        RECT 0.691 0 0.709 0.018 ;
        RECT 0.799 0 0.817 0.018 ;
        RECT 0.907 0 0.925 0.018 ;
        RECT 1.015 0 1.033 0.018 ;
        RECT 1.123 0 1.141 0.018 ;
        RECT 1.1965 0 1.2145 0.018 ;
        RECT 1.557 0 1.575 0.018 ;
        RECT 1.968 0 1.986 0.018 ;
        RECT 2.0705 0 2.0885 0.018 ;
        RECT 2.137 0 2.155 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 2.16 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 2.16 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.193 0.27 1.211 0.288 ;
        RECT 1.5535 0.27 1.5715 0.288 ;
        RECT 1.9615 0.27 1.9795 0.288 ;
        RECT 2.0635 0.27 2.0815 0.288 ;
        RECT 2.137 0.27 2.155 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.128 1.602 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 1.602 0.232 ;
        RECT 1.584 0.125 1.602 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 1.584 0.126 1.602 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 1.584 0.13 1.602 0.148 ;
      LAYER V2 ;
        RECT 1.584 0.135 1.602 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.128 1.224 0.158 ;
        RECT 0.45 0.132 0.468 0.162 ;
      LAYER M2 ;
        RECT 0.45 0.178 1.224 0.196 ;
        RECT 1.206 0.125 1.224 0.196 ;
        RECT 0.45 0.134 0.468 0.196 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.139 0.468 0.157 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.185 1.98 0.203 ;
        RECT 1.962 0.085 1.98 0.203 ;
        RECT 1.233 0.085 1.98 0.103 ;
      LAYER M2 ;
        RECT 1.962 0.125 1.98 0.158 ;
      LAYER M3 ;
        RECT 1.962 0.126 1.98 0.158 ;
      LAYER V1 ;
        RECT 1.962 0.13 1.98 0.148 ;
      LAYER V2 ;
        RECT 1.962 0.135 1.98 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.229 0.765 0.247 ;
      RECT 0.018 0.0865 0.036 0.247 ;
      RECT 0.828 0.0865 0.846 0.15 ;
      RECT 0.018 0.0865 0.846 0.1045 ;
      RECT 0.855 0.042 1.953 0.06 ;
      RECT 1.233 0.228 1.899 0.246 ;
      RECT 0.099 0.042 0.765 0.06 ;
  END
END XNOR2_7x

MACRO XOR2_1x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_1x 0 0 ;
  SIZE 0.54 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.54 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.54 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.0775 0 0.0955 0.018 ;
        RECT 0.187 0 0.205 0.018 ;
        RECT 0.2245 0 0.2425 0.018 ;
        RECT 0.261 0 0.279 0.018 ;
        RECT 0.297 0 0.315 0.018 ;
        RECT 0.348 0 0.366 0.018 ;
        RECT 0.4505 0 0.4685 0.018 ;
        RECT 0.517 0 0.535 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.54 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.041 0.27 0.059 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.113 0.27 0.131 0.288 ;
        RECT 0.149 0.27 0.167 0.288 ;
        RECT 0.185 0.27 0.203 0.288 ;
        RECT 0.221 0.27 0.239 0.288 ;
        RECT 0.2575 0.27 0.2755 0.288 ;
        RECT 0.2935 0.27 0.3115 0.288 ;
        RECT 0.3415 0.27 0.3595 0.288 ;
        RECT 0.4435 0.27 0.4615 0.288 ;
        RECT 0.517 0.27 0.535 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.128 0.252 0.158 ;
        RECT 0.126 0.132 0.144 0.162 ;
      LAYER M2 ;
        RECT 0.126 0.178 0.252 0.196 ;
        RECT 0.234 0.125 0.252 0.196 ;
        RECT 0.126 0.134 0.144 0.196 ;
      LAYER M3 ;
        RECT 0.234 0.126 0.252 0.158 ;
      LAYER V1 ;
        RECT 0.126 0.139 0.144 0.157 ;
        RECT 0.234 0.13 0.252 0.148 ;
      LAYER V2 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.128 0.306 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 0.306 0.232 ;
        RECT 0.288 0.125 0.306 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 0.288 0.126 0.306 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 0.288 0.13 0.306 0.148 ;
      LAYER V2 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.183 0.36 0.201 ;
        RECT 0.342 0.037 0.36 0.201 ;
        RECT 0.207 0.037 0.36 0.055 ;
      LAYER M2 ;
        RECT 0.342 0.125 0.36 0.158 ;
      LAYER M3 ;
        RECT 0.342 0.126 0.36 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.13 0.36 0.148 ;
      LAYER V2 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.233 0.063 0.251 ;
      RECT 0.018 0.087 0.036 0.251 ;
      RECT 0.18 0.087 0.198 0.15 ;
      RECT 0.018 0.087 0.198 0.105 ;
      RECT 0.207 0.226 0.333 0.244 ;
  END
END XOR2_1x

MACRO XOR2_2x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_2x 0 0 ;
  SIZE 0.972 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.972 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.972 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0955 0 0.1135 0.018 ;
        RECT 0.1535 0 0.1715 0.018 ;
        RECT 0.2035 0 0.2215 0.018 ;
        RECT 0.4545 0 0.4725 0.018 ;
        RECT 0.531 0 0.549 0.018 ;
        RECT 0.834 0 0.852 0.018 ;
        RECT 0.8825 0 0.9005 0.018 ;
        RECT 0.949 0 0.967 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 0.972 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 0.972 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.16 0.27 0.178 0.288 ;
        RECT 0.203 0.27 0.221 0.288 ;
        RECT 0.419 0.27 0.437 0.288 ;
        RECT 0.5275 0.27 0.5455 0.288 ;
        RECT 0.72 0.27 0.738 0.288 ;
        RECT 0.8275 0.27 0.8455 0.288 ;
        RECT 0.8755 0.27 0.8935 0.288 ;
        RECT 0.949 0.27 0.967 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.128 0.522 0.158 ;
        RECT 0.18 0.132 0.198 0.162 ;
      LAYER M2 ;
        RECT 0.18 0.178 0.522 0.196 ;
        RECT 0.504 0.125 0.522 0.196 ;
        RECT 0.18 0.134 0.198 0.196 ;
      LAYER M3 ;
        RECT 0.504 0.126 0.522 0.158 ;
      LAYER V1 ;
        RECT 0.18 0.139 0.198 0.157 ;
        RECT 0.504 0.13 0.522 0.148 ;
      LAYER V2 ;
        RECT 0.504 0.135 0.522 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.128 0.738 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 0.738 0.232 ;
        RECT 0.72 0.125 0.738 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.531 0.183 0.846 0.201 ;
        RECT 0.828 0.083 0.846 0.201 ;
        RECT 0.369 0.083 0.846 0.101 ;
      LAYER M2 ;
        RECT 0.828 0.125 0.846 0.158 ;
      LAYER M3 ;
        RECT 0.828 0.126 0.846 0.158 ;
      LAYER V1 ;
        RECT 0.828 0.13 0.846 0.148 ;
      LAYER V2 ;
        RECT 0.828 0.135 0.846 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.19 0.414 0.208 ;
      RECT 0.396 0.132 0.414 0.208 ;
      RECT 0.018 0.087 0.036 0.208 ;
      RECT 0.018 0.087 0.279 0.105 ;
      RECT 0.531 0.04 0.819 0.058 ;
      RECT 0.369 0.233 0.819 0.251 ;
      RECT 0.045 0.233 0.279 0.251 ;
  END
END XOR2_2x

MACRO XOR2_3x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_3x 0 0 ;
  SIZE 1.08 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.08 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.08 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2075 0 0.2255 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.585 0 0.603 0.018 ;
        RECT 0.888 0 0.906 0.018 ;
        RECT 0.9905 0 1.0085 0.018 ;
        RECT 1.057 0 1.075 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.08 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.214 0.27 0.232 0.288 ;
        RECT 0.257 0.27 0.275 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.5815 0.27 0.5995 0.288 ;
        RECT 0.72 0.27 0.738 0.288 ;
        RECT 0.8815 0.27 0.8995 0.288 ;
        RECT 0.9835 0.27 1.0015 0.288 ;
        RECT 1.057 0.27 1.075 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.128 0.576 0.158 ;
        RECT 0.234 0.132 0.252 0.162 ;
      LAYER M2 ;
        RECT 0.234 0.178 0.576 0.196 ;
        RECT 0.558 0.125 0.576 0.196 ;
        RECT 0.234 0.134 0.252 0.196 ;
      LAYER M3 ;
        RECT 0.558 0.126 0.576 0.158 ;
      LAYER V1 ;
        RECT 0.234 0.139 0.252 0.157 ;
        RECT 0.558 0.13 0.576 0.148 ;
      LAYER V2 ;
        RECT 0.558 0.135 0.576 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.128 0.738 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 0.738 0.232 ;
        RECT 0.72 0.125 0.738 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 0.72 0.126 0.738 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 0.72 0.13 0.738 0.148 ;
      LAYER V2 ;
        RECT 0.72 0.135 0.738 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.585 0.183 0.9 0.201 ;
        RECT 0.882 0.083 0.9 0.201 ;
        RECT 0.423 0.083 0.9 0.101 ;
      LAYER M2 ;
        RECT 0.882 0.125 0.9 0.158 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.19 0.414 0.208 ;
      RECT 0.396 0.132 0.414 0.208 ;
      RECT 0.018 0.087 0.036 0.208 ;
      RECT 0.018 0.087 0.333 0.105 ;
      RECT 0.423 0.233 0.873 0.251 ;
      RECT 0.585 0.04 0.819 0.058 ;
      RECT 0.099 0.233 0.333 0.251 ;
  END
END XOR2_3x

MACRO XOR2_5x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_5x 0 0 ;
  SIZE 1.62 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1.62 0.018 ;
      LAYER M2 ;
        RECT 0 0 1.62 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.3155 0 0.3335 0.018 ;
        RECT 0.3655 0 0.3835 0.018 ;
        RECT 0.4735 0 0.4915 0.018 ;
        RECT 0.909 0 0.927 0.018 ;
        RECT 1.428 0 1.446 0.018 ;
        RECT 1.5305 0 1.5485 0.018 ;
        RECT 1.597 0 1.615 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 1.62 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 1.62 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.322 0.27 0.34 0.288 ;
        RECT 0.365 0.27 0.383 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.9055 0.27 0.9235 0.288 ;
        RECT 1.152 0.27 1.17 0.288 ;
        RECT 1.4215 0.27 1.4395 0.288 ;
        RECT 1.5235 0.27 1.5415 0.288 ;
        RECT 1.597 0.27 1.615 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.882 0.128 0.9 0.158 ;
        RECT 0.342 0.132 0.36 0.162 ;
      LAYER M2 ;
        RECT 0.342 0.178 0.9 0.196 ;
        RECT 0.882 0.125 0.9 0.196 ;
        RECT 0.342 0.134 0.36 0.196 ;
      LAYER M3 ;
        RECT 0.882 0.126 0.9 0.158 ;
      LAYER V1 ;
        RECT 0.342 0.139 0.36 0.157 ;
        RECT 0.882 0.13 0.9 0.148 ;
      LAYER V2 ;
        RECT 0.882 0.135 0.9 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.128 1.17 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 1.17 0.232 ;
        RECT 1.152 0.125 1.17 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 1.152 0.126 1.17 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 1.152 0.13 1.17 0.148 ;
      LAYER V2 ;
        RECT 1.152 0.135 1.17 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.909 0.183 1.44 0.201 ;
        RECT 1.422 0.083 1.44 0.201 ;
        RECT 0.639 0.083 1.44 0.101 ;
      LAYER M2 ;
        RECT 1.422 0.125 1.44 0.158 ;
      LAYER M3 ;
        RECT 1.422 0.126 1.44 0.158 ;
      LAYER V1 ;
        RECT 1.422 0.13 1.44 0.148 ;
      LAYER V2 ;
        RECT 1.422 0.135 1.44 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.19 0.63 0.208 ;
      RECT 0.612 0.132 0.63 0.208 ;
      RECT 0.018 0.087 0.036 0.208 ;
      RECT 0.018 0.087 0.549 0.105 ;
      RECT 0.639 0.233 1.413 0.251 ;
      RECT 0.909 0.04 1.359 0.058 ;
      RECT 0.099 0.233 0.549 0.251 ;
  END
END XOR2_5x

MACRO XOR2_7x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_7x 0 0 ;
  SIZE 2.16 BY 0.288 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 2.16 0.018 ;
      LAYER M2 ;
        RECT 0 0 2.16 0.018 ;
      LAYER V1 ;
        RECT 0.005 0 0.023 0.018 ;
        RECT 0.0415 0 0.0595 0.018 ;
        RECT 0.1495 0 0.1675 0.018 ;
        RECT 0.2575 0 0.2755 0.018 ;
        RECT 0.3655 0 0.3835 0.018 ;
        RECT 0.4235 0 0.4415 0.018 ;
        RECT 0.4735 0 0.4915 0.018 ;
        RECT 0.5815 0 0.5995 0.018 ;
        RECT 0.6895 0 0.7075 0.018 ;
        RECT 1.233 0 1.251 0.018 ;
        RECT 1.968 0 1.986 0.018 ;
        RECT 2.0705 0 2.0885 0.018 ;
        RECT 2.137 0 2.155 0.018 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.27 2.16 0.288 ;
      LAYER M2 ;
        RECT 0 0.27 2.16 0.288 ;
      LAYER V1 ;
        RECT 0.005 0.27 0.023 0.288 ;
        RECT 0.077 0.27 0.095 0.288 ;
        RECT 0.43 0.27 0.448 0.288 ;
        RECT 0.473 0.27 0.491 0.288 ;
        RECT 0.581 0.27 0.599 0.288 ;
        RECT 0.689 0.27 0.707 0.288 ;
        RECT 0.797 0.27 0.815 0.288 ;
        RECT 0.905 0.27 0.923 0.288 ;
        RECT 1.013 0.27 1.031 0.288 ;
        RECT 1.121 0.27 1.139 0.288 ;
        RECT 1.2295 0.27 1.2475 0.288 ;
        RECT 1.584 0.27 1.602 0.288 ;
        RECT 1.9615 0.27 1.9795 0.288 ;
        RECT 2.0635 0.27 2.0815 0.288 ;
        RECT 2.137 0.27 2.155 0.288 ;
    END
  END VDD!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.128 1.224 0.158 ;
        RECT 0.45 0.132 0.468 0.162 ;
      LAYER M2 ;
        RECT 0.45 0.178 1.224 0.196 ;
        RECT 1.206 0.125 1.224 0.196 ;
        RECT 0.45 0.134 0.468 0.196 ;
      LAYER M3 ;
        RECT 1.206 0.126 1.224 0.158 ;
      LAYER V1 ;
        RECT 0.45 0.139 0.468 0.157 ;
        RECT 1.206 0.13 1.224 0.148 ;
      LAYER V2 ;
        RECT 1.206 0.135 1.224 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.128 1.602 0.158 ;
        RECT 0.072 0.132 0.09 0.162 ;
      LAYER M2 ;
        RECT 0.072 0.214 1.602 0.232 ;
        RECT 1.584 0.125 1.602 0.232 ;
        RECT 0.072 0.134 0.09 0.232 ;
      LAYER M3 ;
        RECT 1.584 0.126 1.602 0.158 ;
      LAYER V1 ;
        RECT 0.072 0.139 0.09 0.157 ;
        RECT 1.584 0.13 1.602 0.148 ;
      LAYER V2 ;
        RECT 1.584 0.135 1.602 0.153 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.233 0.183 1.98 0.201 ;
        RECT 1.962 0.083 1.98 0.201 ;
        RECT 0.855 0.083 1.98 0.101 ;
      LAYER M2 ;
        RECT 1.962 0.125 1.98 0.158 ;
      LAYER M3 ;
        RECT 1.962 0.126 1.98 0.158 ;
      LAYER V1 ;
        RECT 1.962 0.13 1.98 0.148 ;
      LAYER V2 ;
        RECT 1.962 0.135 1.98 0.153 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 0.018 0.19 0.846 0.208 ;
      RECT 0.828 0.132 0.846 0.208 ;
      RECT 0.018 0.087 0.036 0.208 ;
      RECT 0.018 0.087 0.765 0.105 ;
      RECT 0.855 0.233 1.953 0.251 ;
      RECT 1.233 0.04 1.899 0.058 ;
      RECT 0.099 0.233 0.765 0.251 ;
  END
END XOR2_7x

END LIBRARY
