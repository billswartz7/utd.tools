/Users/bill/version1/utdtools/pgms/cometFlow/tests/test1/riscv/osu035.lef