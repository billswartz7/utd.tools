../../riscv.ckt