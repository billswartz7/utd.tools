/Users/bill/version1/utdtools/pgms/cometFlow/tests/test2/riscv/ASAP7.lef